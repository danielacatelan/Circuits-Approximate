library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

entity M_Mult_AMA3_64 is
 port(
  A    : in std_logic_vector(63 downto 0);
  B    : in std_logic_vector(63 downto 0);
  R    : out std_logic_vector(127 downto 0)
 );
end M_Mult_AMA3_64;

architecture Mult64 of M_Mult_AMA3_64 is

 COMPONENT Soma_AMA3_1
 PORT(
  A : IN std_logic;
  B : IN std_logic;
  Cin : IN std_logic;          
  Cout : OUT std_logic;
  S : OUT std_logic
  );
 END COMPONENT;

 COMPONENT Somador_Exato_1
 PORT(
  A : IN std_logic;
  B : IN std_logic;
  Cin : IN std_logic;          
  Cout : OUT std_logic;
  S : OUT std_logic
  );
 END COMPONENT;
 
signal C : STD_LOGIC_VECTOR (4096 downto 0); --saida das AND
signal Carry : STD_LOGIC_VECTOR (4031 downto 0); -- saida Cout dos somadores
signal E : STD_LOGIC_VECTOR (3906 downto 0); -- Saida S dos somadores

begin
  --b0---
  C(0) <= A(0)and B(0);
  R(0) <= C(0);
  C(1) <= A(1)and B(0); 
  C(2) <= A(2)and B(0);
  C(3) <= A(3)and B(0);
  C(4) <= A(4)and B(0);
  C(5) <= A(5)and B(0);
  C(6) <= A(6)and B(0);
  C(7) <= A(7)and B(0);
  C(8) <= A(8)and B(0);
  C(9) <= A(9)and B(0); 
  C(10) <= A(10)and B(0);
  C(11) <= A(11)and B(0);
  C(12) <= A(12)and B(0);
  C(13) <= A(13)and B(0);
  C(14) <= A(14)and B(0);
  C(15) <= A(15)and B(0);
  C(16) <= A(16)and B(0);
  C(17) <= A(17)and B(0); 
  C(18) <= A(18)and B(0);
  C(19) <= A(19)and B(0);
  C(20) <= A(20)and B(0);
  C(21) <= A(21)and B(0);
  C(22) <= A(22)and B(0);
  C(23) <= A(23)and B(0);
  C(24) <= A(24)and B(0);
  C(25) <= A(25)and B(0); 
  C(26) <= A(26)and B(0);
  C(27) <= A(27)and B(0);
  C(28) <= A(28)and B(0);
  C(29) <= A(29)and B(0);
  C(30) <= A(30)and B(0);
  C(31) <= A(31)and B(0);
  C(32) <= A(32)and B(0);
  C(33) <= A(33)and B(0); 
  C(34) <= A(34)and B(0);
  C(35) <= A(35)and B(0);
  C(36) <= A(36)and B(0);
  C(37) <= A(37)and B(0);
  C(38) <= A(38)and B(0);
  C(39) <= A(39)and B(0);
  C(40) <= A(40)and B(0);
  C(41) <= A(41)and B(0); 
  C(42) <= A(42)and B(0);
  C(43) <= A(43)and B(0);
  C(44) <= A(44)and B(0);
  C(45) <= A(45)and B(0);
  C(46) <= A(46)and B(0);
  C(47) <= A(47)and B(0);  
  C(48) <= A(48)and B(0);
  C(49) <= A(49)and B(0); 
  C(50) <= A(50)and B(0);
  C(51) <= A(51)and B(0);
  C(52) <= A(52)and B(0);
  C(53) <= A(53)and B(0);
  C(54) <= A(54)and B(0);
  C(55) <= A(55)and B(0);
  C(56) <= A(56)and B(0);
  C(57) <= A(57)and B(0); 
  C(58) <= A(58)and B(0);
  C(59) <= A(59)and B(0);
  C(60) <= A(60)and B(0);
  C(61) <= A(61)and B(0);
  C(62) <= A(62)and B(0);
  C(63) <= A(63)and B(0);  
 --b1---
  C(64) <= A(0)and B(1);
  C(65) <= A(1)and B(1); 
  C(66) <= A(2)and B(1);
  C(67) <= A(3)and B(1);
  C(68) <= A(4)and B(1);
  C(69) <= A(5)and B(1);
  C(70) <= A(6)and B(1);
  C(71) <= A(7)and B(1);
  C(72) <= A(8)and B(1);
  C(73) <= A(9)and B(1); 
  C(74) <= A(10)and B(1);
  C(75) <= A(11)and B(1);
  C(76) <= A(12)and B(1);
  C(77) <= A(13)and B(1);
  C(78) <= A(14)and B(1);
  C(79) <= A(15)and B(1);
  C(80) <= A(16)and B(1);
  C(81) <= A(17)and B(1); 
  C(82) <= A(18)and B(1);
  C(83) <= A(19)and B(1);
  C(84) <= A(20)and B(1);
  C(85) <= A(21)and B(1);
  C(86) <= A(22)and B(1);
  C(87) <= A(23)and B(1);
  C(88) <= A(24)and B(1);
  C(89) <= A(25)and B(1); 
  C(90) <= A(26)and B(1);
  C(91) <= A(27)and B(1);
  C(92) <= A(28)and B(1);
  C(93) <= A(29)and B(1);
  C(94) <= A(30)and B(1);
  C(95) <= A(31)and B(1);
  C(96) <= A(32)and B(1);
  C(97) <= A(33)and B(1); 
  C(98) <= A(34)and B(1);
  C(99) <= A(35)and B(1);
  C(100) <= A(36)and B(1);
  C(101) <= A(37)and B(1);
  C(102) <= A(38)and B(1);
  C(103) <= A(39)and B(1);
  C(104) <= A(40)and B(1);
  C(105) <= A(41)and B(1); 
  C(106) <= A(42)and B(1);
  C(107) <= A(43)and B(1);
  C(108) <= A(44)and B(1);
  C(109) <= A(45)and B(1);
  C(110) <= A(46)and B(1);
  C(111) <= A(47)and B(1);  
  C(112) <= A(48)and B(1);
  C(113) <= A(49)and B(1); 
  C(114) <= A(50)and B(1);
  C(115) <= A(51)and B(1);
  C(116) <= A(52)and B(1);
  C(117) <= A(53)and B(1);
  C(118) <= A(54)and B(1);
  C(119) <= A(55)and B(1);
  C(120) <= A(56)and B(1);
  C(121) <= A(57)and B(1); 
  C(122) <= A(58)and B(1);
  C(123) <= A(59)and B(1);
  C(124) <= A(60)and B(1);
  C(125) <= A(61)and B(1);
  C(126) <= A(62)and B(1);
  C(127) <= A(63)and B(1); 
--b2---
  C(128) <= A(0)and B(2);
  C(129) <= A(1)and B(2); 
  C(130) <= A(2)and B(2);
  C(131) <= A(3)and B(2);
  C(132) <= A(4)and B(2);
  C(133) <= A(5)and B(2);
  C(134) <= A(6)and B(2);
  C(135) <= A(7)and B(2);
  C(136) <= A(8)and B(2);
  C(137) <= A(9)and B(2); 
  C(138) <= A(10)and B(2);
  C(139) <= A(11)and B(2);
  C(140) <= A(12)and B(2);
  C(141) <= A(13)and B(2);
  C(142) <= A(14)and B(2);
  C(143) <= A(15)and B(2);
  C(144) <= A(16)and B(2);
  C(145) <= A(17)and B(2); 
  C(146) <= A(18)and B(2);
  C(147) <= A(19)and B(2);
  C(148) <= A(20)and B(2);
  C(149) <= A(21)and B(2);
  C(150) <= A(22)and B(2);
  C(151) <= A(23)and B(2);
  C(152) <= A(24)and B(2);
  C(153) <= A(25)and B(2); 
  C(154) <= A(26)and B(2);
  C(155) <= A(27)and B(2);
  C(156) <= A(28)and B(2);
  C(157) <= A(29)and B(2);
  C(158) <= A(30)and B(2);
  C(159) <= A(31)and B(2);
  C(160) <= A(32)and B(2);
  C(161) <= A(33)and B(2); 
  C(162) <= A(34)and B(2);
  C(163) <= A(35)and B(2);
  C(164) <= A(36)and B(2);
  C(165) <= A(37)and B(2);
  C(166) <= A(38)and B(2);
  C(167) <= A(39)and B(2);
  C(168) <= A(40)and B(2);
  C(169) <= A(41)and B(2); 
  C(170) <= A(42)and B(2);
  C(171) <= A(43)and B(2);
  C(172) <= A(44)and B(2);
  C(173) <= A(45)and B(2);
  C(174) <= A(46)and B(2);
  C(175) <= A(47)and B(2);  
  C(176) <= A(48)and B(2);
  C(177) <= A(49)and B(2); 
  C(178) <= A(50)and B(2);
  C(179) <= A(51)and B(2);
  C(180) <= A(52)and B(2);
  C(181) <= A(53)and B(2);
  C(182) <= A(54)and B(2);
  C(183) <= A(55)and B(2);
  C(184) <= A(56)and B(2);
  C(185) <= A(57)and B(2); 
  C(186) <= A(58)and B(2);
  C(187) <= A(59)and B(2);
  C(188) <= A(60)and B(2);
  C(189) <= A(61)and B(2);
  C(190) <= A(62)and B(2);
  C(191) <= A(63)and B(2);
--b3---
  C(192) <= A(0)and B(3);
  C(193) <= A(1)and B(3); 
  C(194) <= A(2)and B(3);
  C(195) <= A(3)and B(3);
  C(196) <= A(4)and B(3);
  C(197) <= A(5)and B(3);
  C(198) <= A(6)and B(3);
  C(199) <= A(7)and B(3);
  C(200) <= A(8)and B(3);
  C(201) <= A(9)and B(3); 
  C(202) <= A(10)and B(3);
  C(203) <= A(11)and B(3);
  C(204) <= A(12)and B(3);
  C(205) <= A(13)and B(3);
  C(206) <= A(14)and B(3);
  C(207) <= A(15)and B(3);
  C(208) <= A(16)and B(3);
  C(209) <= A(17)and B(3); 
  C(210) <= A(18)and B(3);
  C(211) <= A(19)and B(3);
  C(212) <= A(20)and B(3);
  C(213) <= A(21)and B(3);
  C(214) <= A(22)and B(3);
  C(215) <= A(23)and B(3);
  C(216) <= A(24)and B(3);
  C(217) <= A(25)and B(3); 
  C(218) <= A(26)and B(3);
  C(219) <= A(27)and B(3);
  C(220) <= A(28)and B(3);
  C(221) <= A(29)and B(3);
  C(222) <= A(30)and B(3);
  C(223) <= A(31)and B(3);
  C(224) <= A(32)and B(3);
  C(225) <= A(33)and B(3); 
  C(226) <= A(34)and B(3);
  C(227) <= A(35)and B(3);
  C(228) <= A(36)and B(3);
  C(229) <= A(37)and B(3);
  C(230) <= A(38)and B(3);
  C(231) <= A(39)and B(3);
  C(232) <= A(40)and B(3);
  C(233) <= A(41)and B(3); 
  C(234) <= A(42)and B(3);
  C(235) <= A(43)and B(3);
  C(236) <= A(44)and B(3);
  C(237) <= A(45)and B(3);
  C(238) <= A(46)and B(3);
  C(239) <= A(47)and B(3);  
  C(240) <= A(48)and B(3);
  C(241) <= A(49)and B(3); 
  C(242) <= A(50)and B(3);
  C(243) <= A(51)and B(3);
  C(244) <= A(52)and B(3);
  C(245) <= A(53)and B(3);
  C(246) <= A(54)and B(3);
  C(247) <= A(55)and B(3);
  C(248) <= A(56)and B(3);
  C(249) <= A(57)and B(3); 
  C(250) <= A(58)and B(3);
  C(251) <= A(59)and B(3);
  C(252) <= A(60)and B(3);
  C(253) <= A(61)and B(3);
  C(254) <= A(62)and B(3);
  C(255) <= A(63)and B(3);
--b4---
  C(256) <= A(0)and B(4);
  C(257) <= A(1)and B(4); 
  C(258) <= A(2)and B(4);
  C(259) <= A(3)and B(4);
  C(260) <= A(4)and B(4);
  C(261) <= A(5)and B(4);
  C(262) <= A(6)and B(4);
  C(263) <= A(7)and B(4);
  C(264) <= A(8)and B(4);
  C(265) <= A(9)and B(4); 
  C(266) <= A(10)and B(4);
  C(267) <= A(11)and B(4);
  C(268) <= A(12)and B(4);
  C(269) <= A(13)and B(4);
  C(270) <= A(14)and B(4);
  C(271) <= A(15)and B(4);
  C(272) <= A(16)and B(4);
  C(273) <= A(17)and B(4); 
  C(274) <= A(18)and B(4);
  C(275) <= A(19)and B(4);
  C(276) <= A(20)and B(4);
  C(277) <= A(21)and B(4);
  C(278) <= A(22)and B(4);
  C(279) <= A(23)and B(4);
  C(280) <= A(24)and B(4);
  C(281) <= A(25)and B(4); 
  C(282) <= A(26)and B(4);
  C(283) <= A(27)and B(4);
  C(284) <= A(28)and B(4);
  C(285) <= A(29)and B(4);
  C(286) <= A(30)and B(4);
  C(287) <= A(31)and B(4);
  C(288) <= A(32)and B(4);
  C(289) <= A(33)and B(4); 
  C(290) <= A(34)and B(4);
  C(291) <= A(35)and B(4);
  C(292) <= A(36)and B(4);
  C(293) <= A(37)and B(4);
  C(294) <= A(38)and B(4);
  C(295) <= A(39)and B(4);
  C(296) <= A(40)and B(4);
  C(297) <= A(41)and B(4); 
  C(298) <= A(42)and B(4);
  C(299) <= A(43)and B(4);
  C(300) <= A(44)and B(4);
  C(301) <= A(45)and B(4);
  C(302) <= A(46)and B(4);
  C(303) <= A(47)and B(4);  
  C(304) <= A(48)and B(4);
  C(305) <= A(49)and B(4); 
  C(306) <= A(50)and B(4);
  C(307) <= A(51)and B(4);
  C(308) <= A(52)and B(4);
  C(309) <= A(53)and B(4);
  C(310) <= A(54)and B(4);
  C(311) <= A(55)and B(4);
  C(312) <= A(56)and B(4);
  C(313) <= A(57)and B(4); 
  C(314) <= A(58)and B(4);
  C(315) <= A(59)and B(4);
  C(316) <= A(60)and B(4);
  C(317) <= A(61)and B(4);
  C(318) <= A(62)and B(4);
  C(319) <= A(63)and B(4);
 --b5---
  C(320) <= A(0)and B(5);
  C(321) <= A(1)and B(5); 
  C(322) <= A(2)and B(5);
  C(323) <= A(3)and B(5);
  C(324) <= A(4)and B(5);
  C(325) <= A(5)and B(5);
  C(326) <= A(6)and B(5);
  C(327) <= A(7)and B(5);
  C(328) <= A(8)and B(5);
  C(329) <= A(9)and B(5); 
  C(330) <= A(10)and B(5);
  C(331) <= A(11)and B(5);
  C(332) <= A(12)and B(5);
  C(333) <= A(13)and B(5);
  C(334) <= A(14)and B(5);
  C(335) <= A(15)and B(5);
  C(336) <= A(16)and B(5);
  C(337) <= A(17)and B(5); 
  C(338) <= A(18)and B(5);
  C(339) <= A(19)and B(5);
  C(340) <= A(20)and B(5);
  C(341) <= A(21)and B(5);
  C(342) <= A(22)and B(5);
  C(343) <= A(23)and B(5);
  C(344) <= A(24)and B(5);
  C(345) <= A(25)and B(5); 
  C(346) <= A(26)and B(5);
  C(347) <= A(27)and B(5);
  C(348) <= A(28)and B(5);
  C(349) <= A(29)and B(5);
  C(350) <= A(30)and B(5);
  C(351) <= A(31)and B(5);
  C(352) <= A(32)and B(5);
  C(353) <= A(33)and B(5); 
  C(354) <= A(34)and B(5);
  C(355) <= A(35)and B(5);
  C(356) <= A(36)and B(5);
  C(357) <= A(37)and B(5);
  C(358) <= A(38)and B(5);
  C(359) <= A(39)and B(5);
  C(360) <= A(40)and B(5);
  C(361) <= A(41)and B(5); 
  C(362) <= A(42)and B(5);
  C(363) <= A(43)and B(5);
  C(364) <= A(44)and B(5);
  C(365) <= A(45)and B(5);
  C(366) <= A(46)and B(5);
  C(367) <= A(47)and B(5);  
  C(368) <= A(48)and B(5);
  C(369) <= A(49)and B(5); 
  C(370) <= A(50)and B(5);
  C(371) <= A(51)and B(5);
  C(372) <= A(52)and B(5);
  C(373) <= A(53)and B(5);
  C(374) <= A(54)and B(5);
  C(375) <= A(55)and B(5);
  C(376) <= A(56)and B(5);
  C(377) <= A(57)and B(5); 
  C(378) <= A(58)and B(5);
  C(379) <= A(59)and B(5);
  C(380) <= A(60)and B(5);
  C(381) <= A(61)and B(5);
  C(382) <= A(62)and B(5);
  C(383) <= A(63)and B(5); 
--b6---
  C(384) <= A(0)and B(6);
  C(385) <= A(1)and B(6); 
  C(386) <= A(2)and B(6);
  C(387) <= A(3)and B(6);
  C(388) <= A(4)and B(6);
  C(389) <= A(5)and B(6);
  C(390) <= A(6)and B(6);
  C(391) <= A(7)and B(6);
  C(392) <= A(8)and B(6);
  C(393) <= A(9)and B(6); 
  C(394) <= A(10)and B(6);
  C(395) <= A(11)and B(6);
  C(396) <= A(12)and B(6);
  C(397) <= A(13)and B(6);
  C(398) <= A(14)and B(6);
  C(399) <= A(15)and B(6);
  C(400) <= A(16)and B(6);
  C(401) <= A(17)and B(6); 
  C(402) <= A(18)and B(6);
  C(403) <= A(19)and B(6);
  C(404) <= A(20)and B(6);
  C(405) <= A(21)and B(6);
  C(406) <= A(22)and B(6);
  C(407) <= A(23)and B(6);
  C(408) <= A(24)and B(6);
  C(409) <= A(25)and B(6); 
  C(410) <= A(26)and B(6);
  C(411) <= A(27)and B(6);
  C(412) <= A(28)and B(6);
  C(413) <= A(29)and B(6);
  C(414) <= A(30)and B(6);
  C(415) <= A(31)and B(6);
  C(416) <= A(32)and B(6);
  C(417) <= A(33)and B(6); 
  C(418) <= A(34)and B(6);
  C(419) <= A(35)and B(6);
  C(420) <= A(36)and B(6);
  C(421) <= A(37)and B(6);
  C(422) <= A(38)and B(6);
  C(423) <= A(39)and B(6);
  C(424) <= A(40)and B(6);
  C(425) <= A(41)and B(6); 
  C(426) <= A(42)and B(6);
  C(427) <= A(43)and B(6);
  C(428) <= A(44)and B(6);
  C(429) <= A(45)and B(6);
  C(430) <= A(46)and B(6);
  C(431) <= A(47)and B(6);  
  C(432) <= A(48)and B(6);
  C(433) <= A(49)and B(6); 
  C(434) <= A(50)and B(6);
  C(435) <= A(51)and B(6);
  C(436) <= A(52)and B(6);
  C(437) <= A(53)and B(6);
  C(438) <= A(54)and B(6);
  C(439) <= A(55)and B(6);
  C(440) <= A(56)and B(6);
  C(441) <= A(57)and B(6); 
  C(442) <= A(58)and B(6);
  C(443) <= A(59)and B(6);
  C(444) <= A(60)and B(6);
  C(445) <= A(61)and B(6);
  C(446) <= A(62)and B(6);
  C(447) <= A(63)and B(6);
--b7---
  C(448) <= A(0)and B(7);
  C(449) <= A(1)and B(7); 
  C(450) <= A(2)and B(7);
  C(451) <= A(3)and B(7);
  C(452) <= A(4)and B(7);
  C(453) <= A(5)and B(7);
  C(454) <= A(6)and B(7);
  C(455) <= A(7)and B(7);
  C(456) <= A(8)and B(7);
  C(457) <= A(9)and B(7); 
  C(458) <= A(10)and B(7);
  C(459) <= A(11)and B(7);
  C(460) <= A(12)and B(7);
  C(461) <= A(13)and B(7);
  C(462) <= A(14)and B(7);
  C(463) <= A(15)and B(7);
  C(464) <= A(16)and B(7);
  C(465) <= A(17)and B(7); 
  C(466) <= A(18)and B(7);
  C(467) <= A(19)and B(7);
  C(468) <= A(20)and B(7);
  C(469) <= A(21)and B(7);
  C(470) <= A(22)and B(7);
  C(471) <= A(23)and B(7);
  C(472) <= A(24)and B(7);
  C(473) <= A(25)and B(7); 
  C(474) <= A(26)and B(7);
  C(475) <= A(27)and B(7);
  C(476) <= A(28)and B(7);
  C(477) <= A(29)and B(7);
  C(478) <= A(30)and B(7);
  C(479) <= A(31)and B(7);
  C(480) <= A(32)and B(7);
  C(481) <= A(33)and B(7); 
  C(482) <= A(34)and B(7);
  C(483) <= A(35)and B(7);
  C(484) <= A(36)and B(7);
  C(485) <= A(37)and B(7);
  C(486) <= A(38)and B(7);
  C(487) <= A(39)and B(7);
  C(488) <= A(40)and B(7);
  C(489) <= A(41)and B(7); 
  C(490) <= A(42)and B(7);
  C(491) <= A(43)and B(7);
  C(492) <= A(44)and B(7);
  C(493) <= A(45)and B(7);
  C(494) <= A(46)and B(7);
  C(495) <= A(47)and B(7);  
  C(496) <= A(48)and B(7);
  C(497) <= A(49)and B(7); 
  C(498) <= A(50)and B(7);
  C(499) <= A(51)and B(7);
  C(500) <= A(52)and B(7);
  C(501) <= A(53)and B(7);
  C(502) <= A(54)and B(7);
  C(503) <= A(55)and B(7);
  C(504) <= A(56)and B(7);
  C(505) <= A(57)and B(7); 
  C(506) <= A(58)and B(7);
  C(507) <= A(59)and B(7);
  C(508) <= A(60)and B(7);
  C(509) <= A(61)and B(7);
  C(510) <= A(62)and B(7);
  C(511) <= A(63)and B(7);
--b8---
  C(512) <= A(0)and B(8);
  C(513) <= A(1)and B(8); 
  C(514) <= A(2)and B(8);
  C(515) <= A(3)and B(8);
  C(516) <= A(4)and B(8);
  C(517) <= A(5)and B(8);
  C(518) <= A(6)and B(8);
  C(519) <= A(7)and B(8);
  C(520) <= A(8)and B(8);
  C(521) <= A(9)and B(8); 
  C(522) <= A(10)and B(8);
  C(523) <= A(11)and B(8);
  C(524) <= A(12)and B(8);
  C(525) <= A(13)and B(8);
  C(526) <= A(14)and B(8);
  C(527) <= A(15)and B(8);
  C(528) <= A(16)and B(8);
  C(529) <= A(17)and B(8); 
  C(530) <= A(18)and B(8);
  C(531) <= A(19)and B(8);
  C(532) <= A(20)and B(8);
  C(533) <= A(21)and B(8);
  C(534) <= A(22)and B(8);
  C(535) <= A(23)and B(8);
  C(536) <= A(24)and B(8);
  C(537) <= A(25)and B(8); 
  C(538) <= A(26)and B(8);
  C(539) <= A(27)and B(8);
  C(540) <= A(28)and B(8);
  C(541) <= A(29)and B(8);
  C(542) <= A(30)and B(8);
  C(543) <= A(31)and B(8);
  C(544) <= A(32)and B(8);
  C(545) <= A(33)and B(8); 
  C(546) <= A(34)and B(8);
  C(547) <= A(35)and B(8);
  C(548) <= A(36)and B(8);
  C(549) <= A(37)and B(8);
  C(550) <= A(38)and B(8);
  C(551) <= A(39)and B(8);
  C(552) <= A(40)and B(8);
  C(553) <= A(41)and B(8); 
  C(554) <= A(42)and B(8);
  C(555) <= A(43)and B(8);
  C(556) <= A(44)and B(8);
  C(557) <= A(45)and B(8);
  C(558) <= A(46)and B(8);
  C(559) <= A(47)and B(8);  
  C(560) <= A(48)and B(8);
  C(561) <= A(49)and B(8); 
  C(562) <= A(50)and B(8);
  C(563) <= A(51)and B(8);
  C(564) <= A(52)and B(8);
  C(565) <= A(53)and B(8);
  C(566) <= A(54)and B(8);
  C(567) <= A(55)and B(8);
  C(568) <= A(56)and B(8);
  C(569) <= A(57)and B(8); 
  C(570) <= A(58)and B(8);
  C(571) <= A(59)and B(8);
  C(572) <= A(60)and B(8);
  C(573) <= A(61)and B(8);
  C(574) <= A(62)and B(8);
  C(575) <= A(63)and B(8);
   --b9---
  C(576) <= A(0)and B(9);
  C(577) <= A(1)and B(9); 
  C(578) <= A(2)and B(9);
  C(579) <= A(3)and B(9);
  C(580) <= A(4)and B(9);
  C(581) <= A(5)and B(9);
  C(582) <= A(6)and B(9);
  C(583) <= A(7)and B(9);
  C(584) <= A(8)and B(9);
  C(585) <= A(9)and B(9); 
  C(586) <= A(10)and B(9);
  C(587) <= A(11)and B(9);
  C(588) <= A(12)and B(9);
  C(589) <= A(13)and B(9);
  C(590) <= A(14)and B(9);
  C(591) <= A(15)and B(9);
  C(592) <= A(16)and B(9);
  C(593) <= A(17)and B(9); 
  C(594) <= A(18)and B(9);
  C(595) <= A(19)and B(9);
  C(596) <= A(20)and B(9);
  C(597) <= A(21)and B(9);
  C(598) <= A(22)and B(9);
  C(599) <= A(23)and B(9);
  C(600) <= A(24)and B(9);
  C(601) <= A(25)and B(9); 
  C(602) <= A(26)and B(9);
  C(603) <= A(27)and B(9);
  C(604) <= A(28)and B(9);
  C(605) <= A(29)and B(9);
  C(606) <= A(30)and B(9);
  C(607) <= A(31)and B(9);
  C(608) <= A(32)and B(9);
  C(609) <= A(33)and B(9); 
  C(610) <= A(34)and B(9);
  C(611) <= A(35)and B(9);
  C(612) <= A(36)and B(9);
  C(613) <= A(37)and B(9);
  C(614) <= A(38)and B(9);
  C(615) <= A(39)and B(9);
  C(616) <= A(40)and B(9);
  C(617) <= A(41)and B(9); 
  C(618) <= A(42)and B(9);
  C(619) <= A(43)and B(9);
  C(620) <= A(44)and B(9);
  C(621) <= A(45)and B(9);
  C(622) <= A(46)and B(9);
  C(623) <= A(47)and B(9);  
  C(624) <= A(48)and B(9);
  C(625) <= A(49)and B(9); 
  C(626) <= A(50)and B(9);
  C(627) <= A(51)and B(9);
  C(628) <= A(52)and B(9);
  C(629) <= A(53)and B(9);
  C(630) <= A(54)and B(9);
  C(631) <= A(55)and B(9);
  C(632) <= A(56)and B(9);
  C(633) <= A(57)and B(9); 
  C(634) <= A(58)and B(9);
  C(635) <= A(59)and B(9);
  C(636) <= A(60)and B(9);
  C(637) <= A(61)and B(9);
  C(638) <= A(62)and B(9);
  C(639) <= A(63)and B(9); 
--b10---
  C(640) <= A(0)and B(10);
  C(641) <= A(1)and B(10); 
  C(642) <= A(2)and B(10);
  C(643) <= A(3)and B(10);
  C(644) <= A(4)and B(10);
  C(645) <= A(5)and B(10);
  C(646) <= A(6)and B(10);
  C(647) <= A(7)and B(10);
  C(648) <= A(8)and B(10);
  C(649) <= A(9)and B(10); 
  C(650) <= A(10)and B(10);
  C(651) <= A(11)and B(10);
  C(652) <= A(12)and B(10);
  C(653) <= A(13)and B(10);
  C(654) <= A(14)and B(10);
  C(655) <= A(15)and B(10);
  C(656) <= A(16)and B(10);
  C(657) <= A(17)and B(10); 
  C(658) <= A(18)and B(10);
  C(659) <= A(19)and B(10);
  C(660) <= A(20)and B(10);
  C(661) <= A(21)and B(10);
  C(662) <= A(22)and B(10);
  C(663) <= A(23)and B(10);
  C(664) <= A(24)and B(10);
  C(665) <= A(25)and B(10); 
  C(666) <= A(26)and B(10);
  C(667) <= A(27)and B(10);
  C(668) <= A(28)and B(10);
  C(669) <= A(29)and B(10);
  C(670) <= A(30)and B(10);
  C(671) <= A(31)and B(10);
  C(672) <= A(32)and B(10);
  C(673) <= A(33)and B(10); 
  C(674) <= A(34)and B(10);
  C(675) <= A(35)and B(10);
  C(676) <= A(36)and B(10);
  C(677) <= A(37)and B(10);
  C(678) <= A(38)and B(10);
  C(679) <= A(39)and B(10);
  C(680) <= A(40)and B(10);
  C(681) <= A(41)and B(10); 
  C(682) <= A(42)and B(10);
  C(683) <= A(43)and B(10);
  C(684) <= A(44)and B(10);
  C(685) <= A(45)and B(10);
  C(686) <= A(46)and B(10);
  C(687) <= A(47)and B(10);  
  C(688) <= A(48)and B(10);
  C(689) <= A(49)and B(10); 
  C(690) <= A(50)and B(10);
  C(691) <= A(51)and B(10);
  C(692) <= A(52)and B(10);
  C(693) <= A(53)and B(10);
  C(694) <= A(54)and B(10);
  C(695) <= A(55)and B(10);
  C(696) <= A(56)and B(10);
  C(697) <= A(57)and B(10); 
  C(698) <= A(58)and B(10);
  C(699) <= A(59)and B(10);
  C(700) <= A(60)and B(10);
  C(701) <= A(61)and B(10);
  C(702) <= A(62)and B(10);
  C(703) <= A(63)and B(10);
--b11---
  C(704) <= A(0)and B(11);
  C(705) <= A(1)and B(11); 
  C(706) <= A(2)and B(11);
  C(707) <= A(3)and B(11);
  C(708) <= A(4)and B(11);
  C(709) <= A(5)and B(11);
  C(710) <= A(6)and B(11);
  C(711) <= A(7)and B(11);
  C(712) <= A(8)and B(11);
  C(713) <= A(9)and B(11); 
  C(714) <= A(10)and B(11);
  C(715) <= A(11)and B(11);
  C(716) <= A(12)and B(11);
  C(717) <= A(13)and B(11);
  C(718) <= A(14)and B(11);
  C(719) <= A(15)and B(11);
  C(720) <= A(16)and B(11);
  C(721) <= A(17)and B(11); 
  C(722) <= A(18)and B(11);
  C(723) <= A(19)and B(11);
  C(724) <= A(20)and B(11);
  C(725) <= A(21)and B(11);
  C(726) <= A(22)and B(11);
  C(727) <= A(23)and B(11);
  C(728) <= A(24)and B(11);
  C(729) <= A(25)and B(11); 
  C(730) <= A(26)and B(11);
  C(731) <= A(27)and B(11);
  C(732) <= A(28)and B(11);
  C(733) <= A(29)and B(11);
  C(734) <= A(30)and B(11);
  C(735) <= A(31)and B(11);
  C(736) <= A(32)and B(11);
  C(737) <= A(33)and B(11); 
  C(738) <= A(34)and B(11);
  C(739) <= A(35)and B(11);
  C(740) <= A(36)and B(11);
  C(741) <= A(37)and B(11);
  C(742) <= A(38)and B(11);
  C(743) <= A(39)and B(11);
  C(744) <= A(40)and B(11);
  C(745) <= A(41)and B(11); 
  C(746) <= A(42)and B(11);
  C(747) <= A(43)and B(11);
  C(748) <= A(44)and B(11);
  C(749) <= A(45)and B(11);
  C(750) <= A(46)and B(11);
  C(751) <= A(47)and B(11);  
  C(752) <= A(48)and B(11);
  C(753) <= A(49)and B(11); 
  C(754) <= A(50)and B(11);
  C(755) <= A(51)and B(11);
  C(756) <= A(52)and B(11);
  C(757) <= A(53)and B(11);
  C(758) <= A(54)and B(11);
  C(759) <= A(55)and B(11);
  C(760) <= A(56)and B(11);
  C(761) <= A(57)and B(11); 
  C(762) <= A(58)and B(11);
  C(763) <= A(59)and B(11);
  C(764) <= A(60)and B(11);
  C(765) <= A(61)and B(11);
  C(766) <= A(62)and B(11);
  C(767) <= A(63)and B(11);
--b12---
  C(768) <= A(0)and B(12);
  C(769) <= A(1)and B(12); 
  C(770) <= A(2)and B(12);
  C(771) <= A(3)and B(12);
  C(772) <= A(4)and B(12);
  C(773) <= A(5)and B(12);
  C(774) <= A(6)and B(12);
  C(775) <= A(7)and B(12);
  C(776) <= A(8)and B(12);
  C(777) <= A(9)and B(12); 
  C(778) <= A(10)and B(12);
  C(779) <= A(11)and B(12);
  C(780) <= A(12)and B(12);
  C(781) <= A(13)and B(12);
  C(782) <= A(14)and B(12);
  C(783) <= A(15)and B(12);
  C(784) <= A(16)and B(12);
  C(785) <= A(17)and B(12); 
  C(786) <= A(18)and B(12);
  C(787) <= A(19)and B(12);
  C(788) <= A(20)and B(12);
  C(789) <= A(21)and B(12);
  C(790) <= A(22)and B(12);
  C(791) <= A(23)and B(12);
  C(792) <= A(24)and B(12);
  C(793) <= A(25)and B(12); 
  C(794) <= A(26)and B(12);
  C(795) <= A(27)and B(12);
  C(796) <= A(28)and B(12);
  C(797) <= A(29)and B(12);
  C(798) <= A(30)and B(12);
  C(799) <= A(31)and B(12);
  C(800) <= A(32)and B(12);
  C(801) <= A(33)and B(12); 
  C(802) <= A(34)and B(12);
  C(803) <= A(35)and B(12);
  C(804) <= A(36)and B(12);
  C(805) <= A(37)and B(12);
  C(806) <= A(38)and B(12);
  C(807) <= A(39)and B(12);
  C(808) <= A(40)and B(12);
  C(809) <= A(41)and B(12); 
  C(810) <= A(42)and B(12);
  C(811) <= A(43)and B(12);
  C(812) <= A(44)and B(12);
  C(813) <= A(45)and B(12);
  C(814) <= A(46)and B(12);
  C(815) <= A(47)and B(12);  
  C(816) <= A(48)and B(12);
  C(817) <= A(49)and B(12); 
  C(818) <= A(50)and B(12);
  C(819) <= A(51)and B(12);
  C(820) <= A(52)and B(12);
  C(821) <= A(53)and B(12);
  C(822) <= A(54)and B(12);
  C(823) <= A(55)and B(12);
  C(824) <= A(56)and B(12);
  C(825) <= A(57)and B(12); 
  C(826) <= A(58)and B(12);
  C(827) <= A(59)and B(12);
  C(828) <= A(60)and B(12);
  C(829) <= A(61)and B(12);
  C(830) <= A(62)and B(12);
  C(831) <= A(63)and B(12);
   --b13---
  C(832) <= A(0)and B(13);
  C(833) <= A(1)and B(13); 
  C(834) <= A(2)and B(13);
  C(835) <= A(3)and B(13);
  C(836) <= A(4)and B(13);
  C(837) <= A(5)and B(13);
  C(838) <= A(6)and B(13);
  C(839) <= A(7)and B(13);
  C(840) <= A(8)and B(13);
  C(841) <= A(9)and B(13); 
  C(842) <= A(10)and B(13);
  C(843) <= A(11)and B(13);
  C(844) <= A(12)and B(13);
  C(845) <= A(13)and B(13);
  C(846) <= A(14)and B(13);
  C(847) <= A(15)and B(13);
  C(848) <= A(16)and B(13);
  C(849) <= A(17)and B(13); 
  C(850) <= A(18)and B(13);
  C(851) <= A(19)and B(13);
  C(852) <= A(20)and B(13);
  C(853) <= A(21)and B(13);
  C(854) <= A(22)and B(13);
  C(855) <= A(23)and B(13);
  C(856) <= A(24)and B(13);
  C(857) <= A(25)and B(13); 
  C(858) <= A(26)and B(13);
  C(859) <= A(27)and B(13);
  C(860) <= A(28)and B(13);
  C(861) <= A(29)and B(13);
  C(862) <= A(30)and B(13);
  C(863) <= A(31)and B(13);
  C(864) <= A(32)and B(13);
  C(865) <= A(33)and B(13); 
  C(866) <= A(34)and B(13);
  C(867) <= A(35)and B(13);
  C(868) <= A(36)and B(13);
  C(869) <= A(37)and B(13);
  C(870) <= A(38)and B(13);
  C(871) <= A(39)and B(13);
  C(872) <= A(40)and B(13);
  C(873) <= A(41)and B(13); 
  C(874) <= A(42)and B(13);
  C(875) <= A(43)and B(13);
  C(876) <= A(44)and B(13);
  C(877) <= A(45)and B(13);
  C(878) <= A(46)and B(13);
  C(879) <= A(47)and B(13);  
  C(880) <= A(48)and B(13);
  C(881) <= A(49)and B(13); 
  C(882) <= A(50)and B(13);
  C(883) <= A(51)and B(13);
  C(884) <= A(52)and B(13);
  C(885) <= A(53)and B(13);
  C(886) <= A(54)and B(13);
  C(887) <= A(55)and B(13);
  C(888) <= A(56)and B(13);
  C(889) <= A(57)and B(13); 
  C(890) <= A(58)and B(13);
  C(891) <= A(59)and B(13);
  C(892) <= A(60)and B(13);
  C(893) <= A(61)and B(13);
  C(894) <= A(62)and B(13);
  C(895) <= A(63)and B(13); 
--b14---
  C(896) <= A(0)and B(14);
  C(897) <= A(1)and B(14); 
  C(898) <= A(2)and B(14);
  C(899) <= A(3)and B(14);
  C(900) <= A(4)and B(14);
  C(901) <= A(5)and B(14);
  C(902) <= A(6)and B(14);
  C(903) <= A(7)and B(14);
  C(904) <= A(8)and B(14);
  C(905) <= A(9)and B(14); 
  C(906) <= A(10)and B(14);
  C(907) <= A(11)and B(14);
  C(908) <= A(12)and B(14);
  C(909) <= A(13)and B(14);
  C(910) <= A(14)and B(14);
  C(911) <= A(15)and B(14);
  C(912) <= A(16)and B(14);
  C(913) <= A(17)and B(14); 
  C(914) <= A(18)and B(14);
  C(915) <= A(19)and B(14);
  C(916) <= A(20)and B(14);
  C(917) <= A(21)and B(14);
  C(918) <= A(22)and B(14);
  C(919) <= A(23)and B(14);
  C(920) <= A(24)and B(14);
  C(921) <= A(25)and B(14); 
  C(922) <= A(26)and B(14);
  C(923) <= A(27)and B(14);
  C(924) <= A(28)and B(14);
  C(925) <= A(29)and B(14);
  C(926) <= A(30)and B(14);
  C(927) <= A(31)and B(14);
  C(928) <= A(32)and B(14);
  C(929) <= A(33)and B(14); 
  C(930) <= A(34)and B(14);
  C(931) <= A(35)and B(14);
  C(932) <= A(36)and B(14);
  C(933) <= A(37)and B(14);
  C(934) <= A(38)and B(14);
  C(935) <= A(39)and B(14);
  C(936) <= A(40)and B(14);
  C(937) <= A(41)and B(14); 
  C(938) <= A(42)and B(14);
  C(939) <= A(43)and B(14);
  C(940) <= A(44)and B(14);
  C(941) <= A(45)and B(14);
  C(942) <= A(46)and B(14);
  C(943) <= A(47)and B(14);  
  C(944) <= A(48)and B(14);
  C(945) <= A(49)and B(14); 
  C(946) <= A(50)and B(14);
  C(947) <= A(51)and B(14);
  C(948) <= A(52)and B(14);
  C(949) <= A(53)and B(14);
  C(950) <= A(54)and B(14);
  C(951) <= A(55)and B(14);
  C(952) <= A(56)and B(14);
  C(953) <= A(57)and B(14); 
  C(954) <= A(58)and B(14);
  C(955) <= A(59)and B(14);
  C(956) <= A(60)and B(14);
  C(957) <= A(61)and B(14);
  C(958) <= A(62)and B(14);
  C(959) <= A(63)and B(14);
--b15---
  C(960) <= A(0)and B(15);
  C(961) <= A(1)and B(15); 
  C(962) <= A(2)and B(15);
  C(963) <= A(3)and B(15);
  C(964) <= A(4)and B(15);
  C(965) <= A(5)and B(15);
  C(966) <= A(6)and B(15);
  C(967) <= A(7)and B(15);
  C(968) <= A(8)and B(15);
  C(969) <= A(9)and B(15); 
  C(970) <= A(10)and B(15);
  C(971) <= A(11)and B(15);
  C(972) <= A(12)and B(15);
  C(973) <= A(13)and B(15);
  C(974) <= A(14)and B(15);
  C(975) <= A(15)and B(15);
  C(976) <= A(16)and B(15);
  C(977) <= A(17)and B(15); 
  C(978) <= A(18)and B(15);
  C(979) <= A(19)and B(15);
  C(980) <= A(20)and B(15);
  C(981) <= A(21)and B(15);
  C(982) <= A(22)and B(15);
  C(983) <= A(23)and B(15);
  C(984) <= A(24)and B(15);
  C(985) <= A(25)and B(15); 
  C(986) <= A(26)and B(15);
  C(987) <= A(27)and B(15);
  C(988) <= A(28)and B(15);
  C(989) <= A(29)and B(15);
  C(990) <= A(30)and B(15);
  C(991) <= A(31)and B(15);
  C(992) <= A(32)and B(15);
  C(993) <= A(33)and B(15); 
  C(994) <= A(34)and B(15);
  C(995) <= A(35)and B(15);
  C(996) <= A(36)and B(15);
  C(997) <= A(37)and B(15);
  C(998) <= A(38)and B(15);
  C(999) <= A(39)and B(15);
  C(1000) <= A(40)and B(15);
  C(1001) <= A(41)and B(15); 
  C(1002) <= A(42)and B(15);
  C(1003) <= A(43)and B(15);
  C(1004) <= A(44)and B(15);
  C(1005) <= A(45)and B(15);
  C(1006) <= A(46)and B(15);
  C(1007) <= A(47)and B(15);  
  C(1008) <= A(48)and B(15);
  C(1009) <= A(49)and B(15); 
  C(1010) <= A(50)and B(15);
  C(1011) <= A(51)and B(15);
  C(1012) <= A(52)and B(15);
  C(1013) <= A(53)and B(15);
  C(1014) <= A(54)and B(15);
  C(1015) <= A(55)and B(15);
  C(1016) <= A(56)and B(15);
  C(1017) <= A(57)and B(15); 
  C(1018) <= A(58)and B(15);
  C(1019) <= A(59)and B(15);
  C(1020) <= A(60)and B(15);
  C(1021) <= A(61)and B(15);
  C(1022) <= A(62)and B(15);
  C(1023) <= A(63)and B(15);
--b16---
  C(1024) <= A(0)and B(16);
  C(1025) <= A(1)and B(16); 
  C(1026) <= A(2)and B(16);
  C(1027) <= A(3)and B(16);
  C(1028) <= A(4)and B(16);
  C(1029) <= A(5)and B(16);
  C(1030) <= A(6)and B(16);
  C(1031) <= A(7)and B(16);
  C(1032) <= A(8)and B(16);
  C(1033) <= A(9)and B(16); 
  C(1034) <= A(10)and B(16);
  C(1035) <= A(11)and B(16);
  C(1036) <= A(12)and B(16);
  C(1037) <= A(13)and B(16);
  C(1038) <= A(14)and B(16);
  C(1039) <= A(15)and B(16);
  C(1040) <= A(16)and B(16);
  C(1041) <= A(17)and B(16); 
  C(1042) <= A(18)and B(16);
  C(1043) <= A(19)and B(16);
  C(1044) <= A(20)and B(16);
  C(1045) <= A(21)and B(16);
  C(1046) <= A(22)and B(16);
  C(1047) <= A(23)and B(16);
  C(1048) <= A(24)and B(16);
  C(1049) <= A(25)and B(16); 
  C(1050) <= A(26)and B(16);
  C(1051) <= A(27)and B(16);
  C(1052) <= A(28)and B(16);
  C(1053) <= A(29)and B(16);
  C(1054) <= A(30)and B(16);
  C(1055) <= A(31)and B(16);
  C(1056) <= A(32)and B(16);
  C(1057) <= A(33)and B(16); 
  C(1058) <= A(34)and B(16);
  C(1059) <= A(35)and B(16);
  C(1060) <= A(36)and B(16);
  C(1061) <= A(37)and B(16);
  C(1062) <= A(38)and B(16);
  C(1063) <= A(39)and B(16);
  C(1064) <= A(40)and B(16);
  C(1065) <= A(41)and B(16); 
  C(1066) <= A(42)and B(16);
  C(1067) <= A(43)and B(16);
  C(1068) <= A(44)and B(16);
  C(1069) <= A(45)and B(16);
  C(1070) <= A(46)and B(16);
  C(1071) <= A(47)and B(16);  
  C(1072) <= A(48)and B(16);
  C(1073) <= A(49)and B(16); 
  C(1074) <= A(50)and B(16);
  C(1075) <= A(51)and B(16);
  C(1076) <= A(52)and B(16);
  C(1077) <= A(53)and B(16);
  C(1078) <= A(54)and B(16);
  C(1079) <= A(55)and B(16);
  C(1080) <= A(56)and B(16);
  C(1081) <= A(57)and B(16); 
  C(1082) <= A(58)and B(16);
  C(1083) <= A(59)and B(16);
  C(1084) <= A(60)and B(16);
  C(1085) <= A(61)and B(16);
  C(1086) <= A(62)and B(16);
  C(1087) <= A(63)and B(16);
  --b17---
	C	(	1088	)	<= A(	0	)and B(	17	);
	C	(	1089	)	<= A(	1	)and B(	17	);
	C	(	1090	)	<= A(	2	)and B(	17	);
	C	(	1091	)	<= A(	3	)and B(	17	);
	C	(	1092	)	<= A(	4	)and B(	17	);
	C	(	1093	)	<= A(	5	)and B(	17	);
	C	(	1094	)	<= A(	6	)and B(	17	);
	C	(	1095	)	<= A(	7	)and B(	17	);
	C	(	1096	)	<= A(	8	)and B(	17	);
	C	(	1097	)	<= A(	9	)and B(	17	);
	C	(	1098	)	<= A(	10	)and B(	17	);
	C	(	1099	)	<= A(	11	)and B(	17	);
	C	(	1100	)	<= A(	12	)and B(	17	);
	C	(	1101	)	<= A(	13	)and B(	17	);
	C	(	1102	)	<= A(	14	)and B(	17	);
	C	(	1103	)	<= A(	15	)and B(	17	);
	C	(	1104	)	<= A(	16	)and B(	17	);
	C	(	1105	)	<= A(	17	)and B(	17	);
	C	(	1106	)	<= A(	18	)and B(	17	);
	C	(	1107	)	<= A(	19	)and B(	17	);
	C	(	1108	)	<= A(	20	)and B(	17	);
	C	(	1109	)	<= A(	21	)and B(	17	);
	C	(	1110	)	<= A(	22	)and B(	17	);
	C	(	1111	)	<= A(	23	)and B(	17	);
	C	(	1112	)	<= A(	24	)and B(	17	);
	C	(	1113	)	<= A(	25	)and B(	17	);
	C	(	1114	)	<= A(	26	)and B(	17	);
	C	(	1115	)	<= A(	27	)and B(	17	);
	C	(	1116	)	<= A(	28	)and B(	17	);
	C	(	1117	)	<= A(	29	)and B(	17	);
	C	(	1118	)	<= A(	30	)and B(	17	);
	C	(	1119	)	<= A(	31	)and B(	17	);
	C	(	1120	)	<= A(	32	)and B(	17	);
	C	(	1121	)	<= A(	33	)and B(	17	);
	C	(	1122	)	<= A(	34	)and B(	17	);
	C	(	1123	)	<= A(	35	)and B(	17	);
	C	(	1124	)	<= A(	36	)and B(	17	);
	C	(	1125	)	<= A(	37	)and B(	17	);
	C	(	1126	)	<= A(	38	)and B(	17	);
	C	(	1127	)	<= A(	39	)and B(	17	);
	C	(	1128	)	<= A(	40	)and B(	17	);
	C	(	1129	)	<= A(	41	)and B(	17	);
	C	(	1130	)	<= A(	42	)and B(	17	);
	C	(	1131	)	<= A(	43	)and B(	17	);
	C	(	1132	)	<= A(	44	)and B(	17	);
	C	(	1133	)	<= A(	45	)and B(	17	);
	C	(	1134	)	<= A(	46	)and B(	17	);
	C	(	1135	)	<= A(	47	)and B(	17	);
	C	(	1136	)	<= A(	48	)and B(	17	);
	C	(	1137	)	<= A(	49	)and B(	17	);
	C	(	1138	)	<= A(	50	)and B(	17	);
	C	(	1139	)	<= A(	51	)and B(	17	);
	C	(	1140	)	<= A(	52	)and B(	17	);
	C	(	1141	)	<= A(	53	)and B(	17	);
	C	(	1142	)	<= A(	54	)and B(	17	);
	C	(	1143	)	<= A(	55	)and B(	17	);
	C	(	1144	)	<= A(	56	)and B(	17	);
	C	(	1145	)	<= A(	57	)and B(	17	);
	C	(	1146	)	<= A(	58	)and B(	17	);
	C	(	1147	)	<= A(	59	)and B(	17	);
	C	(	1148	)	<= A(	60	)and B(	17	);
	C	(	1149	)	<= A(	61	)and B(	17	);
	C	(	1150	)	<= A(	62	)and B(	17	);
	C	(	1151	)	<= A(	63	)and B(	17	);

	C	(	1152	)	<= A(	0	)and B(	18	);
	C	(	1153	)	<= A(	1	)and B(	18	);
	C	(	1154	)	<= A(	2	)and B(	18	);
	C	(	1155	)	<= A(	3	)and B(	18	);
	C	(	1156	)	<= A(	4	)and B(	18	);
	C	(	1157	)	<= A(	5	)and B(	18	);
	C	(	1158	)	<= A(	6	)and B(	18	);
	C	(	1159	)	<= A(	7	)and B(	18	);
	C	(	1160	)	<= A(	8	)and B(	18	);
	C	(	1161	)	<= A(	9	)and B(	18	);
	C	(	1162	)	<= A(	10	)and B(	18	);
	C	(	1163	)	<= A(	11	)and B(	18	);
	C	(	1164	)	<= A(	12	)and B(	18	);
	C	(	1165	)	<= A(	13	)and B(	18	);
	C	(	1166	)	<= A(	14	)and B(	18	);
	C	(	1167	)	<= A(	15	)and B(	18	);
	C	(	1168	)	<= A(	16	)and B(	18	);
	C	(	1169	)	<= A(	17	)and B(	18	);
	C	(	1170	)	<= A(	18	)and B(	18	);
	C	(	1171	)	<= A(	19	)and B(	18	);
	C	(	1172	)	<= A(	20	)and B(	18	);
	C	(	1173	)	<= A(	21	)and B(	18	);
	C	(	1174	)	<= A(	22	)and B(	18	);
	C	(	1175	)	<= A(	23	)and B(	18	);
	C	(	1176	)	<= A(	24	)and B(	18	);
	C	(	1177	)	<= A(	25	)and B(	18	);
	C	(	1178	)	<= A(	26	)and B(	18	);
	C	(	1179	)	<= A(	27	)and B(	18	);
	C	(	1180	)	<= A(	28	)and B(	18	);
	C	(	1181	)	<= A(	29	)and B(	18	);
	C	(	1182	)	<= A(	30	)and B(	18	);
	C	(	1183	)	<= A(	31	)and B(	18	);
	C	(	1184	)	<= A(	32	)and B(	18	);
	C	(	1185	)	<= A(	33	)and B(	18	);
	C	(	1186	)	<= A(	34	)and B(	18	);
	C	(	1187	)	<= A(	35	)and B(	18	);
	C	(	1188	)	<= A(	36	)and B(	18	);
	C	(	1189	)	<= A(	37	)and B(	18	);
	C	(	1190	)	<= A(	38	)and B(	18	);
	C	(	1191	)	<= A(	39	)and B(	18	);
	C	(	1192	)	<= A(	40	)and B(	18	);
	C	(	1193	)	<= A(	41	)and B(	18	);
	C	(	1194	)	<= A(	42	)and B(	18	);
	C	(	1195	)	<= A(	43	)and B(	18	);
	C	(	1196	)	<= A(	44	)and B(	18	);
	C	(	1197	)	<= A(	45	)and B(	18	);
	C	(	1198	)	<= A(	46	)and B(	18	);
	C	(	1199	)	<= A(	47	)and B(	18	);
	C	(	1200	)	<= A(	48	)and B(	18	);
	C	(	1201	)	<= A(	49	)and B(	18	);
	C	(	1202	)	<= A(	50	)and B(	18	);
	C	(	1203	)	<= A(	51	)and B(	18	);
	C	(	1204	)	<= A(	52	)and B(	18	);
	C	(	1205	)	<= A(	53	)and B(	18	);
	C	(	1206	)	<= A(	54	)and B(	18	);
	C	(	1207	)	<= A(	55	)and B(	18	);
	C	(	1208	)	<= A(	56	)and B(	18	);
	C	(	1209	)	<= A(	57	)and B(	18	);
	C	(	1210	)	<= A(	58	)and B(	18	);
	C	(	1211	)	<= A(	59	)and B(	18	);
	C	(	1212	)	<= A(	60	)and B(	18	);
	C	(	1213	)	<= A(	61	)and B(	18	);
	C	(	1214	)	<= A(	62	)and B(	18	);
	C	(	1215	)	<= A(	63	)and B(	18	);

	C	(	1216	)	<= A(	0	)and B(	19	);
	C	(	1217	)	<= A(	1	)and B(	19	);
	C	(	1218	)	<= A(	2	)and B(	19	);
	C	(	1219	)	<= A(	3	)and B(	19	);
	C	(	1220	)	<= A(	4	)and B(	19	);
	C	(	1221	)	<= A(	5	)and B(	19	);
	C	(	1222	)	<= A(	6	)and B(	19	);
	C	(	1223	)	<= A(	7	)and B(	19	);
	C	(	1224	)	<= A(	8	)and B(	19	);
	C	(	1225	)	<= A(	9	)and B(	19	);
	C	(	1226	)	<= A(	10	)and B(	19	);
	C	(	1227	)	<= A(	11	)and B(	19	);
	C	(	1228	)	<= A(	12	)and B(	19	);
	C	(	1229	)	<= A(	13	)and B(	19	);
	C	(	1230	)	<= A(	14	)and B(	19	);
	C	(	1231	)	<= A(	15	)and B(	19	);
	C	(	1232	)	<= A(	16	)and B(	19	);
	C	(	1233	)	<= A(	17	)and B(	19	);
	C	(	1234	)	<= A(	18	)and B(	19	);
	C	(	1235	)	<= A(	19	)and B(	19	);
	C	(	1236	)	<= A(	20	)and B(	19	);
	C	(	1237	)	<= A(	21	)and B(	19	);
	C	(	1238	)	<= A(	22	)and B(	19	);
	C	(	1239	)	<= A(	23	)and B(	19	);
	C	(	1240	)	<= A(	24	)and B(	19	);
	C	(	1241	)	<= A(	25	)and B(	19	);
	C	(	1242	)	<= A(	26	)and B(	19	);
	C	(	1243	)	<= A(	27	)and B(	19	);
	C	(	1244	)	<= A(	28	)and B(	19	);
	C	(	1245	)	<= A(	29	)and B(	19	);
	C	(	1246	)	<= A(	30	)and B(	19	);
	C	(	1247	)	<= A(	31	)and B(	19	);
	C	(	1248	)	<= A(	32	)and B(	19	);
	C	(	1249	)	<= A(	33	)and B(	19	);
	C	(	1250	)	<= A(	34	)and B(	19	);
	C	(	1251	)	<= A(	35	)and B(	19	);
	C	(	1252	)	<= A(	36	)and B(	19	);
	C	(	1253	)	<= A(	37	)and B(	19	);
	C	(	1254	)	<= A(	38	)and B(	19	);
	C	(	1255	)	<= A(	39	)and B(	19	);
	C	(	1256	)	<= A(	40	)and B(	19	);
	C	(	1257	)	<= A(	41	)and B(	19	);
	C	(	1258	)	<= A(	42	)and B(	19	);
	C	(	1259	)	<= A(	43	)and B(	19	);
	C	(	1260	)	<= A(	44	)and B(	19	);
	C	(	1261	)	<= A(	45	)and B(	19	);
	C	(	1262	)	<= A(	46	)and B(	19	);
	C	(	1263	)	<= A(	47	)and B(	19	);
	C	(	1264	)	<= A(	48	)and B(	19	);
	C	(	1265	)	<= A(	49	)and B(	19	);
	C	(	1266	)	<= A(	50	)and B(	19	);
	C	(	1267	)	<= A(	51	)and B(	19	);
	C	(	1268	)	<= A(	52	)and B(	19	);
	C	(	1269	)	<= A(	53	)and B(	19	);
	C	(	1270	)	<= A(	54	)and B(	19	);
	C	(	1271	)	<= A(	55	)and B(	19	);
	C	(	1272	)	<= A(	56	)and B(	19	);
	C	(	1273	)	<= A(	57	)and B(	19	);
	C	(	1274	)	<= A(	58	)and B(	19	);
	C	(	1275	)	<= A(	59	)and B(	19	);
	C	(	1276	)	<= A(	60	)and B(	19	);
	C	(	1277	)	<= A(	61	)and B(	19	);
	C	(	1278	)	<= A(	62	)and B(	19	);
	C	(	1279	)	<= A(	63	)and B(	19	);

	C	(	1280	)	<= A(	0	)and B(	20	);
	C	(	1281	)	<= A(	1	)and B(	20	);
	C	(	1282	)	<= A(	2	)and B(	20	);
	C	(	1283	)	<= A(	3	)and B(	20	);
	C	(	1284	)	<= A(	4	)and B(	20	);
	C	(	1285	)	<= A(	5	)and B(	20	);
	C	(	1286	)	<= A(	6	)and B(	20	);
	C	(	1287	)	<= A(	7	)and B(	20	);
	C	(	1288	)	<= A(	8	)and B(	20	);
	C	(	1289	)	<= A(	9	)and B(	20	);
	C	(	1290	)	<= A(	10	)and B(	20	);
	C	(	1291	)	<= A(	11	)and B(	20	);
	C	(	1292	)	<= A(	12	)and B(	20	);
	C	(	1293	)	<= A(	13	)and B(	20	);
	C	(	1294	)	<= A(	14	)and B(	20	);
	C	(	1295	)	<= A(	15	)and B(	20	);
	C	(	1296	)	<= A(	16	)and B(	20	);
	C	(	1297	)	<= A(	17	)and B(	20	);
	C	(	1298	)	<= A(	18	)and B(	20	);
	C	(	1299	)	<= A(	19	)and B(	20	);
	C	(	1300	)	<= A(	20	)and B(	20	);
	C	(	1301	)	<= A(	21	)and B(	20	);
	C	(	1302	)	<= A(	22	)and B(	20	);
	C	(	1303	)	<= A(	23	)and B(	20	);
	C	(	1304	)	<= A(	24	)and B(	20	);
	C	(	1305	)	<= A(	25	)and B(	20	);
	C	(	1306	)	<= A(	26	)and B(	20	);
	C	(	1307	)	<= A(	27	)and B(	20	);
	C	(	1308	)	<= A(	28	)and B(	20	);
	C	(	1309	)	<= A(	29	)and B(	20	);
	C	(	1310	)	<= A(	30	)and B(	20	);
	C	(	1311	)	<= A(	31	)and B(	20	);
	C	(	1312	)	<= A(	32	)and B(	20	);
	C	(	1313	)	<= A(	33	)and B(	20	);
	C	(	1314	)	<= A(	34	)and B(	20	);
	C	(	1315	)	<= A(	35	)and B(	20	);
	C	(	1316	)	<= A(	36	)and B(	20	);
	C	(	1317	)	<= A(	37	)and B(	20	);
	C	(	1318	)	<= A(	38	)and B(	20	);
	C	(	1319	)	<= A(	39	)and B(	20	);
	C	(	1320	)	<= A(	40	)and B(	20	);
	C	(	1321	)	<= A(	41	)and B(	20	);
	C	(	1322	)	<= A(	42	)and B(	20	);
	C	(	1323	)	<= A(	43	)and B(	20	);
	C	(	1324	)	<= A(	44	)and B(	20	);
	C	(	1325	)	<= A(	45	)and B(	20	);
	C	(	1326	)	<= A(	46	)and B(	20	);
	C	(	1327	)	<= A(	47	)and B(	20	);
	C	(	1328	)	<= A(	48	)and B(	20	);
	C	(	1329	)	<= A(	49	)and B(	20	);
	C	(	1330	)	<= A(	50	)and B(	20	);
	C	(	1331	)	<= A(	51	)and B(	20	);
	C	(	1332	)	<= A(	52	)and B(	20	);
	C	(	1333	)	<= A(	53	)and B(	20	);
	C	(	1334	)	<= A(	54	)and B(	20	);
	C	(	1335	)	<= A(	55	)and B(	20	);
	C	(	1336	)	<= A(	56	)and B(	20	);
	C	(	1337	)	<= A(	57	)and B(	20	);
	C	(	1338	)	<= A(	58	)and B(	20	);
	C	(	1339	)	<= A(	59	)and B(	20	);
	C	(	1340	)	<= A(	60	)and B(	20	);
	C	(	1341	)	<= A(	61	)and B(	20	);
	C	(	1342	)	<= A(	62	)and B(	20	);
	C	(	1343	)	<= A(	63	)and B(	20	);

		C	(	1344	)	<= A(	0	)and B(	21	);
	C	(	1345	)	<= A(	1	)and B(	21	);
	C	(	1346	)	<= A(	2	)and B(	21	);
	C	(	1347	)	<= A(	3	)and B(	21	);
	C	(	1348	)	<= A(	4	)and B(	21	);
	C	(	1349	)	<= A(	5	)and B(	21	);
	C	(	1350	)	<= A(	6	)and B(	21	);
	C	(	1351	)	<= A(	7	)and B(	21	);
	C	(	1352	)	<= A(	8	)and B(	21	);
	C	(	1353	)	<= A(	9	)and B(	21	);
	C	(	1354	)	<= A(	10	)and B(	21	);
	C	(	1355	)	<= A(	11	)and B(	21	);
	C	(	1356	)	<= A(	12	)and B(	21	);
	C	(	1357	)	<= A(	13	)and B(	21	);
	C	(	1358	)	<= A(	14	)and B(	21	);
	C	(	1359	)	<= A(	15	)and B(	21	);
	C	(	1360	)	<= A(	16	)and B(	21	);
	C	(	1361	)	<= A(	17	)and B(	21	);
	C	(	1362	)	<= A(	18	)and B(	21	);
	C	(	1363	)	<= A(	19	)and B(	21	);
	C	(	1364	)	<= A(	20	)and B(	21	);
	C	(	1365	)	<= A(	21	)and B(	21	);
	C	(	1366	)	<= A(	22	)and B(	21	);
	C	(	1367	)	<= A(	23	)and B(	21	);
	C	(	1368	)	<= A(	24	)and B(	21	);
	C	(	1369	)	<= A(	25	)and B(	21	);
	C	(	1370	)	<= A(	26	)and B(	21	);
	C	(	1371	)	<= A(	27	)and B(	21	);
	C	(	1372	)	<= A(	28	)and B(	21	);
	C	(	1373	)	<= A(	29	)and B(	21	);
	C	(	1374	)	<= A(	30	)and B(	21	);
	C	(	1375	)	<= A(	31	)and B(	21	);
	C	(	1376	)	<= A(	32	)and B(	21	);
	C	(	1377	)	<= A(	33	)and B(	21	);
	C	(	1378	)	<= A(	34	)and B(	21	);
	C	(	1379	)	<= A(	35	)and B(	21	);
	C	(	1380	)	<= A(	36	)and B(	21	);
	C	(	1381	)	<= A(	37	)and B(	21	);
	C	(	1382	)	<= A(	38	)and B(	21	);
	C	(	1383	)	<= A(	39	)and B(	21	);
	C	(	1384	)	<= A(	40	)and B(	21	);
	C	(	1385	)	<= A(	41	)and B(	21	);
	C	(	1386	)	<= A(	42	)and B(	21	);
	C	(	1387	)	<= A(	43	)and B(	21	);
	C	(	1388	)	<= A(	44	)and B(	21	);
	C	(	1389	)	<= A(	45	)and B(	21	);
	C	(	1390	)	<= A(	46	)and B(	21	);
	C	(	1391	)	<= A(	47	)and B(	21	);
	C	(	1392	)	<= A(	48	)and B(	21	);
	C	(	1393	)	<= A(	49	)and B(	21	);
	C	(	1394	)	<= A(	50	)and B(	21	);
	C	(	1395	)	<= A(	51	)and B(	21	);
	C	(	1396	)	<= A(	52	)and B(	21	);
	C	(	1397	)	<= A(	53	)and B(	21	);
	C	(	1398	)	<= A(	54	)and B(	21	);
	C	(	1399	)	<= A(	55	)and B(	21	);
	C	(	1400	)	<= A(	56	)and B(	21	);
	C	(	1401	)	<= A(	57	)and B(	21	);
	C	(	1402	)	<= A(	58	)and B(	21	);
	C	(	1403	)	<= A(	59	)and B(	21	);
	C	(	1404	)	<= A(	60	)and B(	21	);
	C	(	1405	)	<= A(	61	)and B(	21	);
	C	(	1406	)	<= A(	62	)and B(	21	);
	C	(	1407	)	<= A(	63	)and B(	21	);

	C	(	1408	)	<= A(	0	)and B(	22	);
	C	(	1409	)	<= A(	1	)and B(	22	);
	C	(	1410	)	<= A(	2	)and B(	22	);
	C	(	1411	)	<= A(	3	)and B(	22	);
	C	(	1412	)	<= A(	4	)and B(	22	);
	C	(	1413	)	<= A(	5	)and B(	22	);
	C	(	1414	)	<= A(	6	)and B(	22	);
	C	(	1415	)	<= A(	7	)and B(	22	);
	C	(	1416	)	<= A(	8	)and B(	22	);
	C	(	1417	)	<= A(	9	)and B(	22	);
	C	(	1418	)	<= A(	10	)and B(	22	);
	C	(	1419	)	<= A(	11	)and B(	22	);
	C	(	1420	)	<= A(	12	)and B(	22	);
	C	(	1421	)	<= A(	13	)and B(	22	);
	C	(	1422	)	<= A(	14	)and B(	22	);
	C	(	1423	)	<= A(	15	)and B(	22	);
	C	(	1424	)	<= A(	16	)and B(	22	);
	C	(	1425	)	<= A(	17	)and B(	22	);
	C	(	1426	)	<= A(	18	)and B(	22	);
	C	(	1427	)	<= A(	19	)and B(	22	);
	C	(	1428	)	<= A(	20	)and B(	22	);
	C	(	1429	)	<= A(	21	)and B(	22	);
	C	(	1430	)	<= A(	22	)and B(	22	);
	C	(	1431	)	<= A(	23	)and B(	22	);
	C	(	1432	)	<= A(	24	)and B(	22	);
	C	(	1433	)	<= A(	25	)and B(	22	);
	C	(	1434	)	<= A(	26	)and B(	22	);
	C	(	1435	)	<= A(	27	)and B(	22	);
	C	(	1436	)	<= A(	28	)and B(	22	);
	C	(	1437	)	<= A(	29	)and B(	22	);
	C	(	1438	)	<= A(	30	)and B(	22	);
	C	(	1439	)	<= A(	31	)and B(	22	);
	C	(	1440	)	<= A(	32	)and B(	22	);
	C	(	1441	)	<= A(	33	)and B(	22	);
	C	(	1442	)	<= A(	34	)and B(	22	);
	C	(	1443	)	<= A(	35	)and B(	22	);
	C	(	1444	)	<= A(	36	)and B(	22	);
	C	(	1445	)	<= A(	37	)and B(	22	);
	C	(	1446	)	<= A(	38	)and B(	22	);
	C	(	1447	)	<= A(	39	)and B(	22	);
	C	(	1448	)	<= A(	40	)and B(	22	);
	C	(	1449	)	<= A(	41	)and B(	22	);
	C	(	1450	)	<= A(	42	)and B(	22	);
	C	(	1451	)	<= A(	43	)and B(	22	);
	C	(	1452	)	<= A(	44	)and B(	22	);
	C	(	1453	)	<= A(	45	)and B(	22	);
	C	(	1454	)	<= A(	46	)and B(	22	);
	C	(	1455	)	<= A(	47	)and B(	22	);
	C	(	1456	)	<= A(	48	)and B(	22	);
	C	(	1457	)	<= A(	49	)and B(	22	);
	C	(	1458	)	<= A(	50	)and B(	22	);
	C	(	1459	)	<= A(	51	)and B(	22	);
	C	(	1460	)	<= A(	52	)and B(	22	);
	C	(	1461	)	<= A(	53	)and B(	22	);
	C	(	1462	)	<= A(	54	)and B(	22	);
	C	(	1463	)	<= A(	55	)and B(	22	);
	C	(	1464	)	<= A(	56	)and B(	22	);
	C	(	1465	)	<= A(	57	)and B(	22	);
	C	(	1466	)	<= A(	58	)and B(	22	);
	C	(	1467	)	<= A(	59	)and B(	22	);
	C	(	1468	)	<= A(	60	)and B(	22	);
	C	(	1469	)	<= A(	61	)and B(	22	);
	C	(	1470	)	<= A(	62	)and B(	22	);
	C	(	1471	)	<= A(	63	)and B(	22	);

	C	(	1472	)	<= A(	0	)and B(	23	);
	C	(	1473	)	<= A(	1	)and B(	23	);
	C	(	1474	)	<= A(	2	)and B(	23	);
	C	(	1475	)	<= A(	3	)and B(	23	);
	C	(	1476	)	<= A(	4	)and B(	23	);
	C	(	1477	)	<= A(	5	)and B(	23	);
	C	(	1478	)	<= A(	6	)and B(	23	);
	C	(	1479	)	<= A(	7	)and B(	23	);
	C	(	1480	)	<= A(	8	)and B(	23	);
	C	(	1481	)	<= A(	9	)and B(	23	);
	C	(	1482	)	<= A(	10	)and B(	23	);
	C	(	1483	)	<= A(	11	)and B(	23	);
	C	(	1484	)	<= A(	12	)and B(	23	);
	C	(	1485	)	<= A(	13	)and B(	23	);
	C	(	1486	)	<= A(	14	)and B(	23	);
	C	(	1487	)	<= A(	15	)and B(	23	);
	C	(	1488	)	<= A(	16	)and B(	23	);
	C	(	1489	)	<= A(	17	)and B(	23	);
	C	(	1490	)	<= A(	18	)and B(	23	);
	C	(	1491	)	<= A(	19	)and B(	23	);
	C	(	1492	)	<= A(	20	)and B(	23	);
	C	(	1493	)	<= A(	21	)and B(	23	);
	C	(	1494	)	<= A(	22	)and B(	23	);
	C	(	1495	)	<= A(	23	)and B(	23	);
	C	(	1496	)	<= A(	24	)and B(	23	);
	C	(	1497	)	<= A(	25	)and B(	23	);
	C	(	1498	)	<= A(	26	)and B(	23	);
	C	(	1499	)	<= A(	27	)and B(	23	);
	C	(	1500	)	<= A(	28	)and B(	23	);
	C	(	1501	)	<= A(	29	)and B(	23	);
	C	(	1502	)	<= A(	30	)and B(	23	);
	C	(	1503	)	<= A(	31	)and B(	23	);
	C	(	1504	)	<= A(	32	)and B(	23	);
	C	(	1505	)	<= A(	33	)and B(	23	);
	C	(	1506	)	<= A(	34	)and B(	23	);
	C	(	1507	)	<= A(	35	)and B(	23	);
	C	(	1508	)	<= A(	36	)and B(	23	);
	C	(	1509	)	<= A(	37	)and B(	23	);
	C	(	1510	)	<= A(	38	)and B(	23	);
	C	(	1511	)	<= A(	39	)and B(	23	);
	C	(	1512	)	<= A(	40	)and B(	23	);
	C	(	1513	)	<= A(	41	)and B(	23	);
	C	(	1514	)	<= A(	42	)and B(	23	);
	C	(	1515	)	<= A(	43	)and B(	23	);
	C	(	1516	)	<= A(	44	)and B(	23	);
	C	(	1517	)	<= A(	45	)and B(	23	);
	C	(	1518	)	<= A(	46	)and B(	23	);
	C	(	1519	)	<= A(	47	)and B(	23	);
	C	(	1520	)	<= A(	48	)and B(	23	);
	C	(	1521	)	<= A(	49	)and B(	23	);
	C	(	1522	)	<= A(	50	)and B(	23	);
	C	(	1523	)	<= A(	51	)and B(	23	);
	C	(	1524	)	<= A(	52	)and B(	23	);
	C	(	1525	)	<= A(	53	)and B(	23	);
	C	(	1526	)	<= A(	54	)and B(	23	);
	C	(	1527	)	<= A(	55	)and B(	23	);
	C	(	1528	)	<= A(	56	)and B(	23	);
	C	(	1529	)	<= A(	57	)and B(	23	);
	C	(	1530	)	<= A(	58	)and B(	23	);
	C	(	1531	)	<= A(	59	)and B(	23	);
	C	(	1532	)	<= A(	60	)and B(	23	);
	C	(	1533	)	<= A(	61	)and B(	23	);
	C	(	1534	)	<= A(	62	)and B(	23	);
	C	(	1535	)	<= A(	63	)and B(	23	);

	C	(	1536	)	<= A(	0	)and B(	24	);
	C	(	1537	)	<= A(	1	)and B(	24	);
	C	(	1538	)	<= A(	2	)and B(	24	);
	C	(	1539	)	<= A(	3	)and B(	24	);
	C	(	1540	)	<= A(	4	)and B(	24	);
	C	(	1541	)	<= A(	5	)and B(	24	);
	C	(	1542	)	<= A(	6	)and B(	24	);
	C	(	1543	)	<= A(	7	)and B(	24	);
	C	(	1544	)	<= A(	8	)and B(	24	);
	C	(	1545	)	<= A(	9	)and B(	24	);
	C	(	1546	)	<= A(	10	)and B(	24	);
	C	(	1547	)	<= A(	11	)and B(	24	);
	C	(	1548	)	<= A(	12	)and B(	24	);
	C	(	1549	)	<= A(	13	)and B(	24	);
	C	(	1550	)	<= A(	14	)and B(	24	);
	C	(	1551	)	<= A(	15	)and B(	24	);
	C	(	1552	)	<= A(	16	)and B(	24	);
	C	(	1553	)	<= A(	17	)and B(	24	);
	C	(	1554	)	<= A(	18	)and B(	24	);
	C	(	1555	)	<= A(	19	)and B(	24	);
	C	(	1556	)	<= A(	20	)and B(	24	);
	C	(	1557	)	<= A(	21	)and B(	24	);
	C	(	1558	)	<= A(	22	)and B(	24	);
	C	(	1559	)	<= A(	23	)and B(	24	);
	C	(	1560	)	<= A(	24	)and B(	24	);
	C	(	1561	)	<= A(	25	)and B(	24	);
	C	(	1562	)	<= A(	26	)and B(	24	);
	C	(	1563	)	<= A(	27	)and B(	24	);
	C	(	1564	)	<= A(	28	)and B(	24	);
	C	(	1565	)	<= A(	29	)and B(	24	);
	C	(	1566	)	<= A(	30	)and B(	24	);
	C	(	1567	)	<= A(	31	)and B(	24	);
	C	(	1568	)	<= A(	32	)and B(	24	);
	C	(	1569	)	<= A(	33	)and B(	24	);
	C	(	1570	)	<= A(	34	)and B(	24	);
	C	(	1571	)	<= A(	35	)and B(	24	);
	C	(	1572	)	<= A(	36	)and B(	24	);
	C	(	1573	)	<= A(	37	)and B(	24	);
	C	(	1574	)	<= A(	38	)and B(	24	);
	C	(	1575	)	<= A(	39	)and B(	24	);
	C	(	1576	)	<= A(	40	)and B(	24	);
	C	(	1577	)	<= A(	41	)and B(	24	);
	C	(	1578	)	<= A(	42	)and B(	24	);
	C	(	1579	)	<= A(	43	)and B(	24	);
	C	(	1580	)	<= A(	44	)and B(	24	);
	C	(	1581	)	<= A(	45	)and B(	24	);
	C	(	1582	)	<= A(	46	)and B(	24	);
	C	(	1583	)	<= A(	47	)and B(	24	);
	C	(	1584	)	<= A(	48	)and B(	24	);
	C	(	1585	)	<= A(	49	)and B(	24	);
	C	(	1586	)	<= A(	50	)and B(	24	);
	C	(	1587	)	<= A(	51	)and B(	24	);
	C	(	1588	)	<= A(	52	)and B(	24	);
	C	(	1589	)	<= A(	53	)and B(	24	);
	C	(	1590	)	<= A(	54	)and B(	24	);
	C	(	1591	)	<= A(	55	)and B(	24	);
	C	(	1592	)	<= A(	56	)and B(	24	);
	C	(	1593	)	<= A(	57	)and B(	24	);
	C	(	1594	)	<= A(	58	)and B(	24	);
	C	(	1595	)	<= A(	59	)and B(	24	);
	C	(	1596	)	<= A(	60	)and B(	24	);
	C	(	1597	)	<= A(	61	)and B(	24	);
	C	(	1598	)	<= A(	62	)and B(	24	);
	C	(	1599	)	<= A(	63	)and B(	24	);

	C	(	1600	)	<= A(	0	)and B(	25	);
	C	(	1601	)	<= A(	1	)and B(	25	);
	C	(	1602	)	<= A(	2	)and B(	25	);
	C	(	1603	)	<= A(	3	)and B(	25	);
	C	(	1604	)	<= A(	4	)and B(	25	);
	C	(	1605	)	<= A(	5	)and B(	25	);
	C	(	1606	)	<= A(	6	)and B(	25	);
	C	(	1607	)	<= A(	7	)and B(	25	);
	C	(	1608	)	<= A(	8	)and B(	25	);
	C	(	1609	)	<= A(	9	)and B(	25	);
	C	(	1610	)	<= A(	10	)and B(	25	);
	C	(	1611	)	<= A(	11	)and B(	25	);
	C	(	1612	)	<= A(	12	)and B(	25	);
	C	(	1613	)	<= A(	13	)and B(	25	);
	C	(	1614	)	<= A(	14	)and B(	25	);
	C	(	1615	)	<= A(	15	)and B(	25	);
	C	(	1616	)	<= A(	16	)and B(	25	);
	C	(	1617	)	<= A(	17	)and B(	25	);
	C	(	1618	)	<= A(	18	)and B(	25	);
	C	(	1619	)	<= A(	19	)and B(	25	);
	C	(	1620	)	<= A(	20	)and B(	25	);
	C	(	1621	)	<= A(	21	)and B(	25	);
	C	(	1622	)	<= A(	22	)and B(	25	);
	C	(	1623	)	<= A(	23	)and B(	25	);
	C	(	1624	)	<= A(	24	)and B(	25	);
	C	(	1625	)	<= A(	25	)and B(	25	);
	C	(	1626	)	<= A(	26	)and B(	25	);
	C	(	1627	)	<= A(	27	)and B(	25	);
	C	(	1628	)	<= A(	28	)and B(	25	);
	C	(	1629	)	<= A(	29	)and B(	25	);
	C	(	1630	)	<= A(	30	)and B(	25	);
	C	(	1631	)	<= A(	31	)and B(	25	);
	C	(	1632	)	<= A(	32	)and B(	25	);
	C	(	1633	)	<= A(	33	)and B(	25	);
	C	(	1634	)	<= A(	34	)and B(	25	);
	C	(	1635	)	<= A(	35	)and B(	25	);
	C	(	1636	)	<= A(	36	)and B(	25	);
	C	(	1637	)	<= A(	37	)and B(	25	);
	C	(	1638	)	<= A(	38	)and B(	25	);
	C	(	1639	)	<= A(	39	)and B(	25	);
	C	(	1640	)	<= A(	40	)and B(	25	);
	C	(	1641	)	<= A(	41	)and B(	25	);
	C	(	1642	)	<= A(	42	)and B(	25	);
	C	(	1643	)	<= A(	43	)and B(	25	);
	C	(	1644	)	<= A(	44	)and B(	25	);
	C	(	1645	)	<= A(	45	)and B(	25	);
	C	(	1646	)	<= A(	46	)and B(	25	);
	C	(	1647	)	<= A(	47	)and B(	25	);
	C	(	1648	)	<= A(	48	)and B(	25	);
	C	(	1649	)	<= A(	49	)and B(	25	);
	C	(	1650	)	<= A(	50	)and B(	25	);
	C	(	1651	)	<= A(	51	)and B(	25	);
	C	(	1652	)	<= A(	52	)and B(	25	);
	C	(	1653	)	<= A(	53	)and B(	25	);
	C	(	1654	)	<= A(	54	)and B(	25	);
	C	(	1655	)	<= A(	55	)and B(	25	);
	C	(	1656	)	<= A(	56	)and B(	25	);
	C	(	1657	)	<= A(	57	)and B(	25	);
	C	(	1658	)	<= A(	58	)and B(	25	);
	C	(	1659	)	<= A(	59	)and B(	25	);
	C	(	1660	)	<= A(	60	)and B(	25	);
	C	(	1661	)	<= A(	61	)and B(	25	);
	C	(	1662	)	<= A(	62	)and B(	25	);
	C	(	1663	)	<= A(	63	)and B(	25	);

	C	(	1664	)	<= A(	0	)and B(	26	);
	C	(	1665	)	<= A(	1	)and B(	26	);
	C	(	1666	)	<= A(	2	)and B(	26	);
	C	(	1667	)	<= A(	3	)and B(	26	);
	C	(	1668	)	<= A(	4	)and B(	26	);
	C	(	1669	)	<= A(	5	)and B(	26	);
	C	(	1670	)	<= A(	6	)and B(	26	);
	C	(	1671	)	<= A(	7	)and B(	26	);
	C	(	1672	)	<= A(	8	)and B(	26	);
	C	(	1673	)	<= A(	9	)and B(	26	);
	C	(	1674	)	<= A(	10	)and B(	26	);
	C	(	1675	)	<= A(	11	)and B(	26	);
	C	(	1676	)	<= A(	12	)and B(	26	);
	C	(	1677	)	<= A(	13	)and B(	26	);
	C	(	1678	)	<= A(	14	)and B(	26	);
	C	(	1679	)	<= A(	15	)and B(	26	);
	C	(	1680	)	<= A(	16	)and B(	26	);
	C	(	1681	)	<= A(	17	)and B(	26	);
	C	(	1682	)	<= A(	18	)and B(	26	);
	C	(	1683	)	<= A(	19	)and B(	26	);
	C	(	1684	)	<= A(	20	)and B(	26	);
	C	(	1685	)	<= A(	21	)and B(	26	);
	C	(	1686	)	<= A(	22	)and B(	26	);
	C	(	1687	)	<= A(	23	)and B(	26	);
	C	(	1688	)	<= A(	24	)and B(	26	);
	C	(	1689	)	<= A(	25	)and B(	26	);
	C	(	1690	)	<= A(	26	)and B(	26	);
	C	(	1691	)	<= A(	27	)and B(	26	);
	C	(	1692	)	<= A(	28	)and B(	26	);
	C	(	1693	)	<= A(	29	)and B(	26	);
	C	(	1694	)	<= A(	30	)and B(	26	);
	C	(	1695	)	<= A(	31	)and B(	26	);
	C	(	1696	)	<= A(	32	)and B(	26	);
	C	(	1697	)	<= A(	33	)and B(	26	);
	C	(	1698	)	<= A(	34	)and B(	26	);
	C	(	1699	)	<= A(	35	)and B(	26	);
	C	(	1700	)	<= A(	36	)and B(	26	);
	C	(	1701	)	<= A(	37	)and B(	26	);
	C	(	1702	)	<= A(	38	)and B(	26	);
	C	(	1703	)	<= A(	39	)and B(	26	);
	C	(	1704	)	<= A(	40	)and B(	26	);
	C	(	1705	)	<= A(	41	)and B(	26	);
	C	(	1706	)	<= A(	42	)and B(	26	);
	C	(	1707	)	<= A(	43	)and B(	26	);
	C	(	1708	)	<= A(	44	)and B(	26	);
	C	(	1709	)	<= A(	45	)and B(	26	);
	C	(	1710	)	<= A(	46	)and B(	26	);
	C	(	1711	)	<= A(	47	)and B(	26	);
	C	(	1712	)	<= A(	48	)and B(	26	);
	C	(	1713	)	<= A(	49	)and B(	26	);
	C	(	1714	)	<= A(	50	)and B(	26	);
	C	(	1715	)	<= A(	51	)and B(	26	);
	C	(	1716	)	<= A(	52	)and B(	26	);
	C	(	1717	)	<= A(	53	)and B(	26	);
	C	(	1718	)	<= A(	54	)and B(	26	);
	C	(	1719	)	<= A(	55	)and B(	26	);
	C	(	1720	)	<= A(	56	)and B(	26	);
	C	(	1721	)	<= A(	57	)and B(	26	);
	C	(	1722	)	<= A(	58	)and B(	26	);
	C	(	1723	)	<= A(	59	)and B(	26	);
	C	(	1724	)	<= A(	60	)and B(	26	);
	C	(	1725	)	<= A(	61	)and B(	26	);
	C	(	1726	)	<= A(	62	)and B(	26	);
	C	(	1727	)	<= A(	63	)and B(	26	);

	C	(	1728	)	<= A(	0	)and B(	27	);
	C	(	1729	)	<= A(	1	)and B(	27	);
	C	(	1730	)	<= A(	2	)and B(	27	);
	C	(	1731	)	<= A(	3	)and B(	27	);
	C	(	1732	)	<= A(	4	)and B(	27	);
	C	(	1733	)	<= A(	5	)and B(	27	);
	C	(	1734	)	<= A(	6	)and B(	27	);
	C	(	1735	)	<= A(	7	)and B(	27	);
	C	(	1736	)	<= A(	8	)and B(	27	);
	C	(	1737	)	<= A(	9	)and B(	27	);
	C	(	1738	)	<= A(	10	)and B(	27	);
	C	(	1739	)	<= A(	11	)and B(	27	);
	C	(	1740	)	<= A(	12	)and B(	27	);
	C	(	1741	)	<= A(	13	)and B(	27	);
	C	(	1742	)	<= A(	14	)and B(	27	);
	C	(	1743	)	<= A(	15	)and B(	27	);
	C	(	1744	)	<= A(	16	)and B(	27	);
	C	(	1745	)	<= A(	17	)and B(	27	);
	C	(	1746	)	<= A(	18	)and B(	27	);
	C	(	1747	)	<= A(	19	)and B(	27	);
	C	(	1748	)	<= A(	20	)and B(	27	);
	C	(	1749	)	<= A(	21	)and B(	27	);
	C	(	1750	)	<= A(	22	)and B(	27	);
	C	(	1751	)	<= A(	23	)and B(	27	);
	C	(	1752	)	<= A(	24	)and B(	27	);
	C	(	1753	)	<= A(	25	)and B(	27	);
	C	(	1754	)	<= A(	26	)and B(	27	);
	C	(	1755	)	<= A(	27	)and B(	27	);
	C	(	1756	)	<= A(	28	)and B(	27	);
	C	(	1757	)	<= A(	29	)and B(	27	);
	C	(	1758	)	<= A(	30	)and B(	27	);
	C	(	1759	)	<= A(	31	)and B(	27	);
	C	(	1760	)	<= A(	32	)and B(	27	);
	C	(	1761	)	<= A(	33	)and B(	27	);
	C	(	1762	)	<= A(	34	)and B(	27	);
	C	(	1763	)	<= A(	35	)and B(	27	);
	C	(	1764	)	<= A(	36	)and B(	27	);
	C	(	1765	)	<= A(	37	)and B(	27	);
	C	(	1766	)	<= A(	38	)and B(	27	);
	C	(	1767	)	<= A(	39	)and B(	27	);
	C	(	1768	)	<= A(	40	)and B(	27	);
	C	(	1769	)	<= A(	41	)and B(	27	);
	C	(	1770	)	<= A(	42	)and B(	27	);
	C	(	1771	)	<= A(	43	)and B(	27	);
	C	(	1772	)	<= A(	44	)and B(	27	);
	C	(	1773	)	<= A(	45	)and B(	27	);
	C	(	1774	)	<= A(	46	)and B(	27	);
	C	(	1775	)	<= A(	47	)and B(	27	);
	C	(	1776	)	<= A(	48	)and B(	27	);
	C	(	1777	)	<= A(	49	)and B(	27	);
	C	(	1778	)	<= A(	50	)and B(	27	);
	C	(	1779	)	<= A(	51	)and B(	27	);
	C	(	1780	)	<= A(	52	)and B(	27	);
	C	(	1781	)	<= A(	53	)and B(	27	);
	C	(	1782	)	<= A(	54	)and B(	27	);
	C	(	1783	)	<= A(	55	)and B(	27	);
	C	(	1784	)	<= A(	56	)and B(	27	);
	C	(	1785	)	<= A(	57	)and B(	27	);
	C	(	1786	)	<= A(	58	)and B(	27	);
	C	(	1787	)	<= A(	59	)and B(	27	);
	C	(	1788	)	<= A(	60	)and B(	27	);
	C	(	1789	)	<= A(	61	)and B(	27	);
	C	(	1790	)	<= A(	62	)and B(	27	);
	C	(	1791	)	<= A(	63	)and B(	27	);

	C	(	1792	)	<= A(	0	)and B(	28	);
	C	(	1793	)	<= A(	1	)and B(	28	);
	C	(	1794	)	<= A(	2	)and B(	28	);
	C	(	1795	)	<= A(	3	)and B(	28	);
	C	(	1796	)	<= A(	4	)and B(	28	);
	C	(	1797	)	<= A(	5	)and B(	28	);
	C	(	1798	)	<= A(	6	)and B(	28	);
	C	(	1799	)	<= A(	7	)and B(	28	);
	C	(	1800	)	<= A(	8	)and B(	28	);
	C	(	1801	)	<= A(	9	)and B(	28	);
	C	(	1802	)	<= A(	10	)and B(	28	);
	C	(	1803	)	<= A(	11	)and B(	28	);
	C	(	1804	)	<= A(	12	)and B(	28	);
	C	(	1805	)	<= A(	13	)and B(	28	);
	C	(	1806	)	<= A(	14	)and B(	28	);
	C	(	1807	)	<= A(	15	)and B(	28	);
	C	(	1808	)	<= A(	16	)and B(	28	);
	C	(	1809	)	<= A(	17	)and B(	28	);
	C	(	1810	)	<= A(	18	)and B(	28	);
	C	(	1811	)	<= A(	19	)and B(	28	);
	C	(	1812	)	<= A(	20	)and B(	28	);
	C	(	1813	)	<= A(	21	)and B(	28	);
	C	(	1814	)	<= A(	22	)and B(	28	);
	C	(	1815	)	<= A(	23	)and B(	28	);
	C	(	1816	)	<= A(	24	)and B(	28	);
	C	(	1817	)	<= A(	25	)and B(	28	);
	C	(	1818	)	<= A(	26	)and B(	28	);
	C	(	1819	)	<= A(	27	)and B(	28	);
	C	(	1820	)	<= A(	28	)and B(	28	);
	C	(	1821	)	<= A(	29	)and B(	28	);
	C	(	1822	)	<= A(	30	)and B(	28	);
	C	(	1823	)	<= A(	31	)and B(	28	);
	C	(	1824	)	<= A(	32	)and B(	28	);
	C	(	1825	)	<= A(	33	)and B(	28	);
	C	(	1826	)	<= A(	34	)and B(	28	);
	C	(	1827	)	<= A(	35	)and B(	28	);
	C	(	1828	)	<= A(	36	)and B(	28	);
	C	(	1829	)	<= A(	37	)and B(	28	);
	C	(	1830	)	<= A(	38	)and B(	28	);
	C	(	1831	)	<= A(	39	)and B(	28	);
	C	(	1832	)	<= A(	40	)and B(	28	);
	C	(	1833	)	<= A(	41	)and B(	28	);
	C	(	1834	)	<= A(	42	)and B(	28	);
	C	(	1835	)	<= A(	43	)and B(	28	);
	C	(	1836	)	<= A(	44	)and B(	28	);
	C	(	1837	)	<= A(	45	)and B(	28	);
	C	(	1838	)	<= A(	46	)and B(	28	);
	C	(	1839	)	<= A(	47	)and B(	28	);
	C	(	1840	)	<= A(	48	)and B(	28	);
	C	(	1841	)	<= A(	49	)and B(	28	);
	C	(	1842	)	<= A(	50	)and B(	28	);
	C	(	1843	)	<= A(	51	)and B(	28	);
	C	(	1844	)	<= A(	52	)and B(	28	);
	C	(	1845	)	<= A(	53	)and B(	28	);
	C	(	1846	)	<= A(	54	)and B(	28	);
	C	(	1847	)	<= A(	55	)and B(	28	);
	C	(	1848	)	<= A(	56	)and B(	28	);
	C	(	1849	)	<= A(	57	)and B(	28	);
	C	(	1850	)	<= A(	58	)and B(	28	);
	C	(	1851	)	<= A(	59	)and B(	28	);
	C	(	1852	)	<= A(	60	)and B(	28	);
	C	(	1853	)	<= A(	61	)and B(	28	);
	C	(	1854	)	<= A(	62	)and B(	28	);
	C	(	1855	)	<= A(	63	)and B(	28	);

	C	(	1856	)	<= A(	0	)and B(	29	);
	C	(	1857	)	<= A(	1	)and B(	29	);
	C	(	1858	)	<= A(	2	)and B(	29	);
	C	(	1859	)	<= A(	3	)and B(	29	);
	C	(	1860	)	<= A(	4	)and B(	29	);
	C	(	1861	)	<= A(	5	)and B(	29	);
	C	(	1862	)	<= A(	6	)and B(	29	);
	C	(	1863	)	<= A(	7	)and B(	29	);
	C	(	1864	)	<= A(	8	)and B(	29	);
	C	(	1865	)	<= A(	9	)and B(	29	);
	C	(	1866	)	<= A(	10	)and B(	29	);
	C	(	1867	)	<= A(	11	)and B(	29	);
	C	(	1868	)	<= A(	12	)and B(	29	);
	C	(	1869	)	<= A(	13	)and B(	29	);
	C	(	1870	)	<= A(	14	)and B(	29	);
	C	(	1871	)	<= A(	15	)and B(	29	);
	C	(	1872	)	<= A(	16	)and B(	29	);
	C	(	1873	)	<= A(	17	)and B(	29	);
	C	(	1874	)	<= A(	18	)and B(	29	);
	C	(	1875	)	<= A(	19	)and B(	29	);
	C	(	1876	)	<= A(	20	)and B(	29	);
	C	(	1877	)	<= A(	21	)and B(	29	);
	C	(	1878	)	<= A(	22	)and B(	29	);
	C	(	1879	)	<= A(	23	)and B(	29	);
	C	(	1880	)	<= A(	24	)and B(	29	);
	C	(	1881	)	<= A(	25	)and B(	29	);
	C	(	1882	)	<= A(	26	)and B(	29	);
	C	(	1883	)	<= A(	27	)and B(	29	);
	C	(	1884	)	<= A(	28	)and B(	29	);
	C	(	1885	)	<= A(	29	)and B(	29	);
	C	(	1886	)	<= A(	30	)and B(	29	);
	C	(	1887	)	<= A(	31	)and B(	29	);
	C	(	1888	)	<= A(	32	)and B(	29	);
	C	(	1889	)	<= A(	33	)and B(	29	);
	C	(	1890	)	<= A(	34	)and B(	29	);
	C	(	1891	)	<= A(	35	)and B(	29	);
	C	(	1892	)	<= A(	36	)and B(	29	);
	C	(	1893	)	<= A(	37	)and B(	29	);
	C	(	1894	)	<= A(	38	)and B(	29	);
	C	(	1895	)	<= A(	39	)and B(	29	);
	C	(	1896	)	<= A(	40	)and B(	29	);
	C	(	1897	)	<= A(	41	)and B(	29	);
	C	(	1898	)	<= A(	42	)and B(	29	);
	C	(	1899	)	<= A(	43	)and B(	29	);
	C	(	1900	)	<= A(	44	)and B(	29	);
	C	(	1901	)	<= A(	45	)and B(	29	);
	C	(	1902	)	<= A(	46	)and B(	29	);
	C	(	1903	)	<= A(	47	)and B(	29	);
	C	(	1904	)	<= A(	48	)and B(	29	);
	C	(	1905	)	<= A(	49	)and B(	29	);
	C	(	1906	)	<= A(	50	)and B(	29	);
	C	(	1907	)	<= A(	51	)and B(	29	);
	C	(	1908	)	<= A(	52	)and B(	29	);
	C	(	1909	)	<= A(	53	)and B(	29	);
	C	(	1910	)	<= A(	54	)and B(	29	);
	C	(	1911	)	<= A(	55	)and B(	29	);
	C	(	1912	)	<= A(	56	)and B(	29	);
	C	(	1913	)	<= A(	57	)and B(	29	);
	C	(	1914	)	<= A(	58	)and B(	29	);
	C	(	1915	)	<= A(	59	)and B(	29	);
	C	(	1916	)	<= A(	60	)and B(	29	);
	C	(	1917	)	<= A(	61	)and B(	29	);
	C	(	1918	)	<= A(	62	)and B(	29	);
	C	(	1919	)	<= A(	63	)and B(	29	);

	C	(	1920	)	<= A(	0	)and B(	30	);
	C	(	1921	)	<= A(	1	)and B(	30	);
	C	(	1922	)	<= A(	2	)and B(	30	);
	C	(	1923	)	<= A(	3	)and B(	30	);
	C	(	1924	)	<= A(	4	)and B(	30	);
	C	(	1925	)	<= A(	5	)and B(	30	);
	C	(	1926	)	<= A(	6	)and B(	30	);
	C	(	1927	)	<= A(	7	)and B(	30	);
	C	(	1928	)	<= A(	8	)and B(	30	);
	C	(	1929	)	<= A(	9	)and B(	30	);
	C	(	1930	)	<= A(	10	)and B(	30	);
	C	(	1931	)	<= A(	11	)and B(	30	);
	C	(	1932	)	<= A(	12	)and B(	30	);
	C	(	1933	)	<= A(	13	)and B(	30	);
	C	(	1934	)	<= A(	14	)and B(	30	);
	C	(	1935	)	<= A(	15	)and B(	30	);
	C	(	1936	)	<= A(	16	)and B(	30	);
	C	(	1937	)	<= A(	17	)and B(	30	);
	C	(	1938	)	<= A(	18	)and B(	30	);
	C	(	1939	)	<= A(	19	)and B(	30	);
	C	(	1940	)	<= A(	20	)and B(	30	);
	C	(	1941	)	<= A(	21	)and B(	30	);
	C	(	1942	)	<= A(	22	)and B(	30	);
	C	(	1943	)	<= A(	23	)and B(	30	);
	C	(	1944	)	<= A(	24	)and B(	30	);
	C	(	1945	)	<= A(	25	)and B(	30	);
	C	(	1946	)	<= A(	26	)and B(	30	);
	C	(	1947	)	<= A(	27	)and B(	30	);
	C	(	1948	)	<= A(	28	)and B(	30	);
	C	(	1949	)	<= A(	29	)and B(	30	);
	C	(	1950	)	<= A(	30	)and B(	30	);
	C	(	1951	)	<= A(	31	)and B(	30	);
	C	(	1952	)	<= A(	32	)and B(	30	);
	C	(	1953	)	<= A(	33	)and B(	30	);
	C	(	1954	)	<= A(	34	)and B(	30	);
	C	(	1955	)	<= A(	35	)and B(	30	);
	C	(	1956	)	<= A(	36	)and B(	30	);
	C	(	1957	)	<= A(	37	)and B(	30	);
	C	(	1958	)	<= A(	38	)and B(	30	);
	C	(	1959	)	<= A(	39	)and B(	30	);
	C	(	1960	)	<= A(	40	)and B(	30	);
	C	(	1961	)	<= A(	41	)and B(	30	);
	C	(	1962	)	<= A(	42	)and B(	30	);
	C	(	1963	)	<= A(	43	)and B(	30	);
	C	(	1964	)	<= A(	44	)and B(	30	);
	C	(	1965	)	<= A(	45	)and B(	30	);
	C	(	1966	)	<= A(	46	)and B(	30	);
	C	(	1967	)	<= A(	47	)and B(	30	);
	C	(	1968	)	<= A(	48	)and B(	30	);
	C	(	1969	)	<= A(	49	)and B(	30	);
	C	(	1970	)	<= A(	50	)and B(	30	);
	C	(	1971	)	<= A(	51	)and B(	30	);
	C	(	1972	)	<= A(	52	)and B(	30	);
	C	(	1973	)	<= A(	53	)and B(	30	);
	C	(	1974	)	<= A(	54	)and B(	30	);
	C	(	1975	)	<= A(	55	)and B(	30	);
	C	(	1976	)	<= A(	56	)and B(	30	);
	C	(	1977	)	<= A(	57	)and B(	30	);
	C	(	1978	)	<= A(	58	)and B(	30	);
	C	(	1979	)	<= A(	59	)and B(	30	);
	C	(	1980	)	<= A(	60	)and B(	30	);
	C	(	1981	)	<= A(	61	)and B(	30	);
	C	(	1982	)	<= A(	62	)and B(	30	);
	C	(	1983	)	<= A(	63	)and B(	30	);

	C	(	1984	)	<= A(	0	)and B(	31	);
	C	(	1985	)	<= A(	1	)and B(	31	);
	C	(	1986	)	<= A(	2	)and B(	31	);
	C	(	1987	)	<= A(	3	)and B(	31	);
	C	(	1988	)	<= A(	4	)and B(	31	);
	C	(	1989	)	<= A(	5	)and B(	31	);
	C	(	1990	)	<= A(	6	)and B(	31	);
	C	(	1991	)	<= A(	7	)and B(	31	);
	C	(	1992	)	<= A(	8	)and B(	31	);
	C	(	1993	)	<= A(	9	)and B(	31	);
	C	(	1994	)	<= A(	10	)and B(	31	);
	C	(	1995	)	<= A(	11	)and B(	31	);
	C	(	1996	)	<= A(	12	)and B(	31	);
	C	(	1997	)	<= A(	13	)and B(	31	);
	C	(	1998	)	<= A(	14	)and B(	31	);
	C	(	1999	)	<= A(	15	)and B(	31	);
	C	(	2000	)	<= A(	16	)and B(	31	);
	C	(	2001	)	<= A(	17	)and B(	31	);
	C	(	2002	)	<= A(	18	)and B(	31	);
	C	(	2003	)	<= A(	19	)and B(	31	);
	C	(	2004	)	<= A(	20	)and B(	31	);
	C	(	2005	)	<= A(	21	)and B(	31	);
	C	(	2006	)	<= A(	22	)and B(	31	);
	C	(	2007	)	<= A(	23	)and B(	31	);
	C	(	2008	)	<= A(	24	)and B(	31	);
	C	(	2009	)	<= A(	25	)and B(	31	);
	C	(	2010	)	<= A(	26	)and B(	31	);
	C	(	2011	)	<= A(	27	)and B(	31	);
	C	(	2012	)	<= A(	28	)and B(	31	);
	C	(	2013	)	<= A(	29	)and B(	31	);
	C	(	2014	)	<= A(	30	)and B(	31	);
	C	(	2015	)	<= A(	31	)and B(	31	);
	C	(	2016	)	<= A(	32	)and B(	31	);
	C	(	2017	)	<= A(	33	)and B(	31	);
	C	(	2018	)	<= A(	34	)and B(	31	);
	C	(	2019	)	<= A(	35	)and B(	31	);
	C	(	2020	)	<= A(	36	)and B(	31	);
	C	(	2021	)	<= A(	37	)and B(	31	);
	C	(	2022	)	<= A(	38	)and B(	31	);
	C	(	2023	)	<= A(	39	)and B(	31	);
	C	(	2024	)	<= A(	40	)and B(	31	);
	C	(	2025	)	<= A(	41	)and B(	31	);
	C	(	2026	)	<= A(	42	)and B(	31	);
	C	(	2027	)	<= A(	43	)and B(	31	);
	C	(	2028	)	<= A(	44	)and B(	31	);
	C	(	2029	)	<= A(	45	)and B(	31	);
	C	(	2030	)	<= A(	46	)and B(	31	);
	C	(	2031	)	<= A(	47	)and B(	31	);
	C	(	2032	)	<= A(	48	)and B(	31	);
	C	(	2033	)	<= A(	49	)and B(	31	);
	C	(	2034	)	<= A(	50	)and B(	31	);
	C	(	2035	)	<= A(	51	)and B(	31	);
	C	(	2036	)	<= A(	52	)and B(	31	);
	C	(	2037	)	<= A(	53	)and B(	31	);
	C	(	2038	)	<= A(	54	)and B(	31	);
	C	(	2039	)	<= A(	55	)and B(	31	);
	C	(	2040	)	<= A(	56	)and B(	31	);
	C	(	2041	)	<= A(	57	)and B(	31	);
	C	(	2042	)	<= A(	58	)and B(	31	);
	C	(	2043	)	<= A(	59	)and B(	31	);
	C	(	2044	)	<= A(	60	)and B(	31	);
	C	(	2045	)	<= A(	61	)and B(	31	);
	C	(	2046	)	<= A(	62	)and B(	31	);
	C	(	2047	)	<= A(	63	)and B(	31	);

	C	(	2048	)	<= A(	0	)and B(	32	);
	C	(	2049	)	<= A(	1	)and B(	32	);
	C	(	2050	)	<= A(	2	)and B(	32	);
	C	(	2051	)	<= A(	3	)and B(	32	);
	C	(	2052	)	<= A(	4	)and B(	32	);
	C	(	2053	)	<= A(	5	)and B(	32	);
	C	(	2054	)	<= A(	6	)and B(	32	);
	C	(	2055	)	<= A(	7	)and B(	32	);
	C	(	2056	)	<= A(	8	)and B(	32	);
	C	(	2057	)	<= A(	9	)and B(	32	);
	C	(	2058	)	<= A(	10	)and B(	32	);
	C	(	2059	)	<= A(	11	)and B(	32	);
	C	(	2060	)	<= A(	12	)and B(	32	);
	C	(	2061	)	<= A(	13	)and B(	32	);
	C	(	2062	)	<= A(	14	)and B(	32	);
	C	(	2063	)	<= A(	15	)and B(	32	);
	C	(	2064	)	<= A(	16	)and B(	32	);
	C	(	2065	)	<= A(	17	)and B(	32	);
	C	(	2066	)	<= A(	18	)and B(	32	);
	C	(	2067	)	<= A(	19	)and B(	32	);
	C	(	2068	)	<= A(	20	)and B(	32	);
	C	(	2069	)	<= A(	21	)and B(	32	);
	C	(	2070	)	<= A(	22	)and B(	32	);
	C	(	2071	)	<= A(	23	)and B(	32	);
	C	(	2072	)	<= A(	24	)and B(	32	);
	C	(	2073	)	<= A(	25	)and B(	32	);
	C	(	2074	)	<= A(	26	)and B(	32	);
	C	(	2075	)	<= A(	27	)and B(	32	);
	C	(	2076	)	<= A(	28	)and B(	32	);
	C	(	2077	)	<= A(	29	)and B(	32	);
	C	(	2078	)	<= A(	30	)and B(	32	);
	C	(	2079	)	<= A(	31	)and B(	32	);
	C	(	2080	)	<= A(	32	)and B(	32	);
	C	(	2081	)	<= A(	33	)and B(	32	);
	C	(	2082	)	<= A(	34	)and B(	32	);
	C	(	2083	)	<= A(	35	)and B(	32	);
	C	(	2084	)	<= A(	36	)and B(	32	);
	C	(	2085	)	<= A(	37	)and B(	32	);
	C	(	2086	)	<= A(	38	)and B(	32	);
	C	(	2087	)	<= A(	39	)and B(	32	);
	C	(	2088	)	<= A(	40	)and B(	32	);
	C	(	2089	)	<= A(	41	)and B(	32	);
	C	(	2090	)	<= A(	42	)and B(	32	);
	C	(	2091	)	<= A(	43	)and B(	32	);
	C	(	2092	)	<= A(	44	)and B(	32	);
	C	(	2093	)	<= A(	45	)and B(	32	);
	C	(	2094	)	<= A(	46	)and B(	32	);
	C	(	2095	)	<= A(	47	)and B(	32	);
	C	(	2096	)	<= A(	48	)and B(	32	);
	C	(	2097	)	<= A(	49	)and B(	32	);
	C	(	2098	)	<= A(	50	)and B(	32	);
	C	(	2099	)	<= A(	51	)and B(	32	);
	C	(	2100	)	<= A(	52	)and B(	32	);
	C	(	2101	)	<= A(	53	)and B(	32	);
	C	(	2102	)	<= A(	54	)and B(	32	);
	C	(	2103	)	<= A(	55	)and B(	32	);
	C	(	2104	)	<= A(	56	)and B(	32	);
	C	(	2105	)	<= A(	57	)and B(	32	);
	C	(	2106	)	<= A(	58	)and B(	32	);
	C	(	2107	)	<= A(	59	)and B(	32	);
	C	(	2108	)	<= A(	60	)and B(	32	);
	C	(	2109	)	<= A(	61	)and B(	32	);
	C	(	2110	)	<= A(	62	)and B(	32	);
	C	(	2111	)	<= A(	63	)and B(	32	);

	C	(	2112	)	<= A(	0	)and B(	33	);
	C	(	2113	)	<= A(	1	)and B(	33	);
	C	(	2114	)	<= A(	2	)and B(	33	);
	C	(	2115	)	<= A(	3	)and B(	33	);
	C	(	2116	)	<= A(	4	)and B(	33	);
	C	(	2117	)	<= A(	5	)and B(	33	);
	C	(	2118	)	<= A(	6	)and B(	33	);
	C	(	2119	)	<= A(	7	)and B(	33	);
	C	(	2120	)	<= A(	8	)and B(	33	);
	C	(	2121	)	<= A(	9	)and B(	33	);
	C	(	2122	)	<= A(	10	)and B(	33	);
	C	(	2123	)	<= A(	11	)and B(	33	);
	C	(	2124	)	<= A(	12	)and B(	33	);
	C	(	2125	)	<= A(	13	)and B(	33	);
	C	(	2126	)	<= A(	14	)and B(	33	);
	C	(	2127	)	<= A(	15	)and B(	33	);
	C	(	2128	)	<= A(	16	)and B(	33	);
	C	(	2129	)	<= A(	17	)and B(	33	);
	C	(	2130	)	<= A(	18	)and B(	33	);
	C	(	2131	)	<= A(	19	)and B(	33	);
	C	(	2132	)	<= A(	20	)and B(	33	);
	C	(	2133	)	<= A(	21	)and B(	33	);
	C	(	2134	)	<= A(	22	)and B(	33	);
	C	(	2135	)	<= A(	23	)and B(	33	);
	C	(	2136	)	<= A(	24	)and B(	33	);
	C	(	2137	)	<= A(	25	)and B(	33	);
	C	(	2138	)	<= A(	26	)and B(	33	);
	C	(	2139	)	<= A(	27	)and B(	33	);
	C	(	2140	)	<= A(	28	)and B(	33	);
	C	(	2141	)	<= A(	29	)and B(	33	);
	C	(	2142	)	<= A(	30	)and B(	33	);
	C	(	2143	)	<= A(	31	)and B(	33	);
	C	(	2144	)	<= A(	32	)and B(	33	);
	C	(	2145	)	<= A(	33	)and B(	33	);
	C	(	2146	)	<= A(	34	)and B(	33	);
	C	(	2147	)	<= A(	35	)and B(	33	);
	C	(	2148	)	<= A(	36	)and B(	33	);
	C	(	2149	)	<= A(	37	)and B(	33	);
	C	(	2150	)	<= A(	38	)and B(	33	);
	C	(	2151	)	<= A(	39	)and B(	33	);
	C	(	2152	)	<= A(	40	)and B(	33	);
	C	(	2153	)	<= A(	41	)and B(	33	);
	C	(	2154	)	<= A(	42	)and B(	33	);
	C	(	2155	)	<= A(	43	)and B(	33	);
	C	(	2156	)	<= A(	44	)and B(	33	);
	C	(	2157	)	<= A(	45	)and B(	33	);
	C	(	2158	)	<= A(	46	)and B(	33	);
	C	(	2159	)	<= A(	47	)and B(	33	);
	C	(	2160	)	<= A(	48	)and B(	33	);
	C	(	2161	)	<= A(	49	)and B(	33	);
	C	(	2162	)	<= A(	50	)and B(	33	);
	C	(	2163	)	<= A(	51	)and B(	33	);
	C	(	2164	)	<= A(	52	)and B(	33	);
	C	(	2165	)	<= A(	53	)and B(	33	);
	C	(	2166	)	<= A(	54	)and B(	33	);
	C	(	2167	)	<= A(	55	)and B(	33	);
	C	(	2168	)	<= A(	56	)and B(	33	);
	C	(	2169	)	<= A(	57	)and B(	33	);
	C	(	2170	)	<= A(	58	)and B(	33	);
	C	(	2171	)	<= A(	59	)and B(	33	);
	C	(	2172	)	<= A(	60	)and B(	33	);
	C	(	2173	)	<= A(	61	)and B(	33	);
	C	(	2174	)	<= A(	62	)and B(	33	);
	C	(	2175	)	<= A(	63	)and B(	33	);

	C	(	2176	)	<= A(	0	)and B(	34	);
	C	(	2177	)	<= A(	1	)and B(	34	);
	C	(	2178	)	<= A(	2	)and B(	34	);
	C	(	2179	)	<= A(	3	)and B(	34	);
	C	(	2180	)	<= A(	4	)and B(	34	);
	C	(	2181	)	<= A(	5	)and B(	34	);
	C	(	2182	)	<= A(	6	)and B(	34	);
	C	(	2183	)	<= A(	7	)and B(	34	);
	C	(	2184	)	<= A(	8	)and B(	34	);
	C	(	2185	)	<= A(	9	)and B(	34	);
	C	(	2186	)	<= A(	10	)and B(	34	);
	C	(	2187	)	<= A(	11	)and B(	34	);
	C	(	2188	)	<= A(	12	)and B(	34	);
	C	(	2189	)	<= A(	13	)and B(	34	);
	C	(	2190	)	<= A(	14	)and B(	34	);
	C	(	2191	)	<= A(	15	)and B(	34	);
	C	(	2192	)	<= A(	16	)and B(	34	);
	C	(	2193	)	<= A(	17	)and B(	34	);
	C	(	2194	)	<= A(	18	)and B(	34	);
	C	(	2195	)	<= A(	19	)and B(	34	);
	C	(	2196	)	<= A(	20	)and B(	34	);
	C	(	2197	)	<= A(	21	)and B(	34	);
	C	(	2198	)	<= A(	22	)and B(	34	);
	C	(	2199	)	<= A(	23	)and B(	34	);
	C	(	2200	)	<= A(	24	)and B(	34	);
	C	(	2201	)	<= A(	25	)and B(	34	);
	C	(	2202	)	<= A(	26	)and B(	34	);
	C	(	2203	)	<= A(	27	)and B(	34	);
	C	(	2204	)	<= A(	28	)and B(	34	);
	C	(	2205	)	<= A(	29	)and B(	34	);
	C	(	2206	)	<= A(	30	)and B(	34	);
	C	(	2207	)	<= A(	31	)and B(	34	);
	C	(	2208	)	<= A(	32	)and B(	34	);
	C	(	2209	)	<= A(	33	)and B(	34	);
	C	(	2210	)	<= A(	34	)and B(	34	);
	C	(	2211	)	<= A(	35	)and B(	34	);
	C	(	2212	)	<= A(	36	)and B(	34	);
	C	(	2213	)	<= A(	37	)and B(	34	);
	C	(	2214	)	<= A(	38	)and B(	34	);
	C	(	2215	)	<= A(	39	)and B(	34	);
	C	(	2216	)	<= A(	40	)and B(	34	);
	C	(	2217	)	<= A(	41	)and B(	34	);
	C	(	2218	)	<= A(	42	)and B(	34	);
	C	(	2219	)	<= A(	43	)and B(	34	);
	C	(	2220	)	<= A(	44	)and B(	34	);
	C	(	2221	)	<= A(	45	)and B(	34	);
	C	(	2222	)	<= A(	46	)and B(	34	);
	C	(	2223	)	<= A(	47	)and B(	34	);
	C	(	2224	)	<= A(	48	)and B(	34	);
	C	(	2225	)	<= A(	49	)and B(	34	);
	C	(	2226	)	<= A(	50	)and B(	34	);
	C	(	2227	)	<= A(	51	)and B(	34	);
	C	(	2228	)	<= A(	52	)and B(	34	);
	C	(	2229	)	<= A(	53	)and B(	34	);
	C	(	2230	)	<= A(	54	)and B(	34	);
	C	(	2231	)	<= A(	55	)and B(	34	);
	C	(	2232	)	<= A(	56	)and B(	34	);
	C	(	2233	)	<= A(	57	)and B(	34	);
	C	(	2234	)	<= A(	58	)and B(	34	);
	C	(	2235	)	<= A(	59	)and B(	34	);
	C	(	2236	)	<= A(	60	)and B(	34	);
	C	(	2237	)	<= A(	61	)and B(	34	);
	C	(	2238	)	<= A(	62	)and B(	34	);
	C	(	2239	)	<= A(	63	)and B(	34	);

	C	(	2240	)	<= A(	0	)and B(	35	);
	C	(	2241	)	<= A(	1	)and B(	35	);
	C	(	2242	)	<= A(	2	)and B(	35	);
	C	(	2243	)	<= A(	3	)and B(	35	);
	C	(	2244	)	<= A(	4	)and B(	35	);
	C	(	2245	)	<= A(	5	)and B(	35	);
	C	(	2246	)	<= A(	6	)and B(	35	);
	C	(	2247	)	<= A(	7	)and B(	35	);
	C	(	2248	)	<= A(	8	)and B(	35	);
	C	(	2249	)	<= A(	9	)and B(	35	);
	C	(	2250	)	<= A(	10	)and B(	35	);
	C	(	2251	)	<= A(	11	)and B(	35	);
	C	(	2252	)	<= A(	12	)and B(	35	);
	C	(	2253	)	<= A(	13	)and B(	35	);
	C	(	2254	)	<= A(	14	)and B(	35	);
	C	(	2255	)	<= A(	15	)and B(	35	);
	C	(	2256	)	<= A(	16	)and B(	35	);
	C	(	2257	)	<= A(	17	)and B(	35	);
	C	(	2258	)	<= A(	18	)and B(	35	);
	C	(	2259	)	<= A(	19	)and B(	35	);
	C	(	2260	)	<= A(	20	)and B(	35	);
	C	(	2261	)	<= A(	21	)and B(	35	);
	C	(	2262	)	<= A(	22	)and B(	35	);
	C	(	2263	)	<= A(	23	)and B(	35	);
	C	(	2264	)	<= A(	24	)and B(	35	);
	C	(	2265	)	<= A(	25	)and B(	35	);
	C	(	2266	)	<= A(	26	)and B(	35	);
	C	(	2267	)	<= A(	27	)and B(	35	);
	C	(	2268	)	<= A(	28	)and B(	35	);
	C	(	2269	)	<= A(	29	)and B(	35	);
	C	(	2270	)	<= A(	30	)and B(	35	);
	C	(	2271	)	<= A(	31	)and B(	35	);
	C	(	2272	)	<= A(	32	)and B(	35	);
	C	(	2273	)	<= A(	33	)and B(	35	);
	C	(	2274	)	<= A(	34	)and B(	35	);
	C	(	2275	)	<= A(	35	)and B(	35	);
	C	(	2276	)	<= A(	36	)and B(	35	);
	C	(	2277	)	<= A(	37	)and B(	35	);
	C	(	2278	)	<= A(	38	)and B(	35	);
	C	(	2279	)	<= A(	39	)and B(	35	);
	C	(	2280	)	<= A(	40	)and B(	35	);
	C	(	2281	)	<= A(	41	)and B(	35	);
	C	(	2282	)	<= A(	42	)and B(	35	);
	C	(	2283	)	<= A(	43	)and B(	35	);
	C	(	2284	)	<= A(	44	)and B(	35	);
	C	(	2285	)	<= A(	45	)and B(	35	);
	C	(	2286	)	<= A(	46	)and B(	35	);
	C	(	2287	)	<= A(	47	)and B(	35	);
	C	(	2288	)	<= A(	48	)and B(	35	);
	C	(	2289	)	<= A(	49	)and B(	35	);
	C	(	2290	)	<= A(	50	)and B(	35	);
	C	(	2291	)	<= A(	51	)and B(	35	);
	C	(	2292	)	<= A(	52	)and B(	35	);
	C	(	2293	)	<= A(	53	)and B(	35	);
	C	(	2294	)	<= A(	54	)and B(	35	);
	C	(	2295	)	<= A(	55	)and B(	35	);
	C	(	2296	)	<= A(	56	)and B(	35	);
	C	(	2297	)	<= A(	57	)and B(	35	);
	C	(	2298	)	<= A(	58	)and B(	35	);
	C	(	2299	)	<= A(	59	)and B(	35	);
	C	(	2300	)	<= A(	60	)and B(	35	);
	C	(	2301	)	<= A(	61	)and B(	35	);
	C	(	2302	)	<= A(	62	)and B(	35	);
	C	(	2303	)	<= A(	63	)and B(	35	);

	C	(	2304	)	<= A(	0	)and B(	36	);
	C	(	2305	)	<= A(	1	)and B(	36	);
	C	(	2306	)	<= A(	2	)and B(	36	);
	C	(	2307	)	<= A(	3	)and B(	36	);
	C	(	2308	)	<= A(	4	)and B(	36	);
	C	(	2309	)	<= A(	5	)and B(	36	);
	C	(	2310	)	<= A(	6	)and B(	36	);
	C	(	2311	)	<= A(	7	)and B(	36	);
	C	(	2312	)	<= A(	8	)and B(	36	);
	C	(	2313	)	<= A(	9	)and B(	36	);
	C	(	2314	)	<= A(	10	)and B(	36	);
	C	(	2315	)	<= A(	11	)and B(	36	);
	C	(	2316	)	<= A(	12	)and B(	36	);
	C	(	2317	)	<= A(	13	)and B(	36	);
	C	(	2318	)	<= A(	14	)and B(	36	);
	C	(	2319	)	<= A(	15	)and B(	36	);
	C	(	2320	)	<= A(	16	)and B(	36	);
	C	(	2321	)	<= A(	17	)and B(	36	);
	C	(	2322	)	<= A(	18	)and B(	36	);
	C	(	2323	)	<= A(	19	)and B(	36	);
	C	(	2324	)	<= A(	20	)and B(	36	);
	C	(	2325	)	<= A(	21	)and B(	36	);
	C	(	2326	)	<= A(	22	)and B(	36	);
	C	(	2327	)	<= A(	23	)and B(	36	);
	C	(	2328	)	<= A(	24	)and B(	36	);
	C	(	2329	)	<= A(	25	)and B(	36	);
	C	(	2330	)	<= A(	26	)and B(	36	);
	C	(	2331	)	<= A(	27	)and B(	36	);
	C	(	2332	)	<= A(	28	)and B(	36	);
	C	(	2333	)	<= A(	29	)and B(	36	);
	C	(	2334	)	<= A(	30	)and B(	36	);
	C	(	2335	)	<= A(	31	)and B(	36	);
	C	(	2336	)	<= A(	32	)and B(	36	);
	C	(	2337	)	<= A(	33	)and B(	36	);
	C	(	2338	)	<= A(	34	)and B(	36	);
	C	(	2339	)	<= A(	35	)and B(	36	);
	C	(	2340	)	<= A(	36	)and B(	36	);
	C	(	2341	)	<= A(	37	)and B(	36	);
	C	(	2342	)	<= A(	38	)and B(	36	);
	C	(	2343	)	<= A(	39	)and B(	36	);
	C	(	2344	)	<= A(	40	)and B(	36	);
	C	(	2345	)	<= A(	41	)and B(	36	);
	C	(	2346	)	<= A(	42	)and B(	36	);
	C	(	2347	)	<= A(	43	)and B(	36	);
	C	(	2348	)	<= A(	44	)and B(	36	);
	C	(	2349	)	<= A(	45	)and B(	36	);
	C	(	2350	)	<= A(	46	)and B(	36	);
	C	(	2351	)	<= A(	47	)and B(	36	);
	C	(	2352	)	<= A(	48	)and B(	36	);
	C	(	2353	)	<= A(	49	)and B(	36	);
	C	(	2354	)	<= A(	50	)and B(	36	);
	C	(	2355	)	<= A(	51	)and B(	36	);
	C	(	2356	)	<= A(	52	)and B(	36	);
	C	(	2357	)	<= A(	53	)and B(	36	);
	C	(	2358	)	<= A(	54	)and B(	36	);
	C	(	2359	)	<= A(	55	)and B(	36	);
	C	(	2360	)	<= A(	56	)and B(	36	);
	C	(	2361	)	<= A(	57	)and B(	36	);
	C	(	2362	)	<= A(	58	)and B(	36	);
	C	(	2363	)	<= A(	59	)and B(	36	);
	C	(	2364	)	<= A(	60	)and B(	36	);
	C	(	2365	)	<= A(	61	)and B(	36	);
	C	(	2366	)	<= A(	62	)and B(	36	);
	C	(	2367	)	<= A(	63	)and B(	36	);

	C	(	2368	)	<= A(	0	)and B(	37	);
	C	(	2369	)	<= A(	1	)and B(	37	);
	C	(	2370	)	<= A(	2	)and B(	37	);
	C	(	2371	)	<= A(	3	)and B(	37	);
	C	(	2372	)	<= A(	4	)and B(	37	);
	C	(	2373	)	<= A(	5	)and B(	37	);
	C	(	2374	)	<= A(	6	)and B(	37	);
	C	(	2375	)	<= A(	7	)and B(	37	);
	C	(	2376	)	<= A(	8	)and B(	37	);
	C	(	2377	)	<= A(	9	)and B(	37	);
	C	(	2378	)	<= A(	10	)and B(	37	);
	C	(	2379	)	<= A(	11	)and B(	37	);
	C	(	2380	)	<= A(	12	)and B(	37	);
	C	(	2381	)	<= A(	13	)and B(	37	);
	C	(	2382	)	<= A(	14	)and B(	37	);
	C	(	2383	)	<= A(	15	)and B(	37	);
	C	(	2384	)	<= A(	16	)and B(	37	);
	C	(	2385	)	<= A(	17	)and B(	37	);
	C	(	2386	)	<= A(	18	)and B(	37	);
	C	(	2387	)	<= A(	19	)and B(	37	);
	C	(	2388	)	<= A(	20	)and B(	37	);
	C	(	2389	)	<= A(	21	)and B(	37	);
	C	(	2390	)	<= A(	22	)and B(	37	);
	C	(	2391	)	<= A(	23	)and B(	37	);
	C	(	2392	)	<= A(	24	)and B(	37	);
	C	(	2393	)	<= A(	25	)and B(	37	);
	C	(	2394	)	<= A(	26	)and B(	37	);
	C	(	2395	)	<= A(	27	)and B(	37	);
	C	(	2396	)	<= A(	28	)and B(	37	);
	C	(	2397	)	<= A(	29	)and B(	37	);
	C	(	2398	)	<= A(	30	)and B(	37	);
	C	(	2399	)	<= A(	31	)and B(	37	);
	C	(	2400	)	<= A(	32	)and B(	37	);
	C	(	2401	)	<= A(	33	)and B(	37	);
	C	(	2402	)	<= A(	34	)and B(	37	);
	C	(	2403	)	<= A(	35	)and B(	37	);
	C	(	2404	)	<= A(	36	)and B(	37	);
	C	(	2405	)	<= A(	37	)and B(	37	);
	C	(	2406	)	<= A(	38	)and B(	37	);
	C	(	2407	)	<= A(	39	)and B(	37	);
	C	(	2408	)	<= A(	40	)and B(	37	);
	C	(	2409	)	<= A(	41	)and B(	37	);
	C	(	2410	)	<= A(	42	)and B(	37	);
	C	(	2411	)	<= A(	43	)and B(	37	);
	C	(	2412	)	<= A(	44	)and B(	37	);
	C	(	2413	)	<= A(	45	)and B(	37	);
	C	(	2414	)	<= A(	46	)and B(	37	);
	C	(	2415	)	<= A(	47	)and B(	37	);
	C	(	2416	)	<= A(	48	)and B(	37	);
	C	(	2417	)	<= A(	49	)and B(	37	);
	C	(	2418	)	<= A(	50	)and B(	37	);
	C	(	2419	)	<= A(	51	)and B(	37	);
	C	(	2420	)	<= A(	52	)and B(	37	);
	C	(	2421	)	<= A(	53	)and B(	37	);
	C	(	2422	)	<= A(	54	)and B(	37	);
	C	(	2423	)	<= A(	55	)and B(	37	);
	C	(	2424	)	<= A(	56	)and B(	37	);
	C	(	2425	)	<= A(	57	)and B(	37	);
	C	(	2426	)	<= A(	58	)and B(	37	);
	C	(	2427	)	<= A(	59	)and B(	37	);
	C	(	2428	)	<= A(	60	)and B(	37	);
	C	(	2429	)	<= A(	61	)and B(	37	);
	C	(	2430	)	<= A(	62	)and B(	37	);
	C	(	2431	)	<= A(	63	)and B(	37	);

	C	(	2432	)	<= A(	0	)and B(	38	);
	C	(	2433	)	<= A(	1	)and B(	38	);
	C	(	2434	)	<= A(	2	)and B(	38	);
	C	(	2435	)	<= A(	3	)and B(	38	);
	C	(	2436	)	<= A(	4	)and B(	38	);
	C	(	2437	)	<= A(	5	)and B(	38	);
	C	(	2438	)	<= A(	6	)and B(	38	);
	C	(	2439	)	<= A(	7	)and B(	38	);
	C	(	2440	)	<= A(	8	)and B(	38	);
	C	(	2441	)	<= A(	9	)and B(	38	);
	C	(	2442	)	<= A(	10	)and B(	38	);
	C	(	2443	)	<= A(	11	)and B(	38	);
	C	(	2444	)	<= A(	12	)and B(	38	);
	C	(	2445	)	<= A(	13	)and B(	38	);
	C	(	2446	)	<= A(	14	)and B(	38	);
	C	(	2447	)	<= A(	15	)and B(	38	);
	C	(	2448	)	<= A(	16	)and B(	38	);
	C	(	2449	)	<= A(	17	)and B(	38	);
	C	(	2450	)	<= A(	18	)and B(	38	);
	C	(	2451	)	<= A(	19	)and B(	38	);
	C	(	2452	)	<= A(	20	)and B(	38	);
	C	(	2453	)	<= A(	21	)and B(	38	);
	C	(	2454	)	<= A(	22	)and B(	38	);
	C	(	2455	)	<= A(	23	)and B(	38	);
	C	(	2456	)	<= A(	24	)and B(	38	);
	C	(	2457	)	<= A(	25	)and B(	38	);
	C	(	2458	)	<= A(	26	)and B(	38	);
	C	(	2459	)	<= A(	27	)and B(	38	);
	C	(	2460	)	<= A(	28	)and B(	38	);
	C	(	2461	)	<= A(	29	)and B(	38	);
	C	(	2462	)	<= A(	30	)and B(	38	);
	C	(	2463	)	<= A(	31	)and B(	38	);
	C	(	2464	)	<= A(	32	)and B(	38	);
	C	(	2465	)	<= A(	33	)and B(	38	);
	C	(	2466	)	<= A(	34	)and B(	38	);
	C	(	2467	)	<= A(	35	)and B(	38	);
	C	(	2468	)	<= A(	36	)and B(	38	);
	C	(	2469	)	<= A(	37	)and B(	38	);
	C	(	2470	)	<= A(	38	)and B(	38	);
	C	(	2471	)	<= A(	39	)and B(	38	);
	C	(	2472	)	<= A(	40	)and B(	38	);
	C	(	2473	)	<= A(	41	)and B(	38	);
	C	(	2474	)	<= A(	42	)and B(	38	);
	C	(	2475	)	<= A(	43	)and B(	38	);
	C	(	2476	)	<= A(	44	)and B(	38	);
	C	(	2477	)	<= A(	45	)and B(	38	);
	C	(	2478	)	<= A(	46	)and B(	38	);
	C	(	2479	)	<= A(	47	)and B(	38	);
	C	(	2480	)	<= A(	48	)and B(	38	);
	C	(	2481	)	<= A(	49	)and B(	38	);
	C	(	2482	)	<= A(	50	)and B(	38	);
	C	(	2483	)	<= A(	51	)and B(	38	);
	C	(	2484	)	<= A(	52	)and B(	38	);
	C	(	2485	)	<= A(	53	)and B(	38	);
	C	(	2486	)	<= A(	54	)and B(	38	);
	C	(	2487	)	<= A(	55	)and B(	38	);
	C	(	2488	)	<= A(	56	)and B(	38	);
	C	(	2489	)	<= A(	57	)and B(	38	);
	C	(	2490	)	<= A(	58	)and B(	38	);
	C	(	2491	)	<= A(	59	)and B(	38	);
	C	(	2492	)	<= A(	60	)and B(	38	);
	C	(	2493	)	<= A(	61	)and B(	38	);
	C	(	2494	)	<= A(	62	)and B(	38	);
	C	(	2495	)	<= A(	63	)and B(	38	);

	C	(	2496	)	<= A(	0	)and B(	39	);
	C	(	2497	)	<= A(	1	)and B(	39	);
	C	(	2498	)	<= A(	2	)and B(	39	);
	C	(	2499	)	<= A(	3	)and B(	39	);
	C	(	2500	)	<= A(	4	)and B(	39	);
	C	(	2501	)	<= A(	5	)and B(	39	);
	C	(	2502	)	<= A(	6	)and B(	39	);
	C	(	2503	)	<= A(	7	)and B(	39	);
	C	(	2504	)	<= A(	8	)and B(	39	);
	C	(	2505	)	<= A(	9	)and B(	39	);
	C	(	2506	)	<= A(	10	)and B(	39	);
	C	(	2507	)	<= A(	11	)and B(	39	);
	C	(	2508	)	<= A(	12	)and B(	39	);
	C	(	2509	)	<= A(	13	)and B(	39	);
	C	(	2510	)	<= A(	14	)and B(	39	);
	C	(	2511	)	<= A(	15	)and B(	39	);
	C	(	2512	)	<= A(	16	)and B(	39	);
	C	(	2513	)	<= A(	17	)and B(	39	);
	C	(	2514	)	<= A(	18	)and B(	39	);
	C	(	2515	)	<= A(	19	)and B(	39	);
	C	(	2516	)	<= A(	20	)and B(	39	);
	C	(	2517	)	<= A(	21	)and B(	39	);
	C	(	2518	)	<= A(	22	)and B(	39	);
	C	(	2519	)	<= A(	23	)and B(	39	);
	C	(	2520	)	<= A(	24	)and B(	39	);
	C	(	2521	)	<= A(	25	)and B(	39	);
	C	(	2522	)	<= A(	26	)and B(	39	);
	C	(	2523	)	<= A(	27	)and B(	39	);
	C	(	2524	)	<= A(	28	)and B(	39	);
	C	(	2525	)	<= A(	29	)and B(	39	);
	C	(	2526	)	<= A(	30	)and B(	39	);
	C	(	2527	)	<= A(	31	)and B(	39	);
	C	(	2528	)	<= A(	32	)and B(	39	);
	C	(	2529	)	<= A(	33	)and B(	39	);
	C	(	2530	)	<= A(	34	)and B(	39	);
	C	(	2531	)	<= A(	35	)and B(	39	);
	C	(	2532	)	<= A(	36	)and B(	39	);
	C	(	2533	)	<= A(	37	)and B(	39	);
	C	(	2534	)	<= A(	38	)and B(	39	);
	C	(	2535	)	<= A(	39	)and B(	39	);
	C	(	2536	)	<= A(	40	)and B(	39	);
	C	(	2537	)	<= A(	41	)and B(	39	);
	C	(	2538	)	<= A(	42	)and B(	39	);
	C	(	2539	)	<= A(	43	)and B(	39	);
	C	(	2540	)	<= A(	44	)and B(	39	);
	C	(	2541	)	<= A(	45	)and B(	39	);
	C	(	2542	)	<= A(	46	)and B(	39	);
	C	(	2543	)	<= A(	47	)and B(	39	);
	C	(	2544	)	<= A(	48	)and B(	39	);
	C	(	2545	)	<= A(	49	)and B(	39	);
	C	(	2546	)	<= A(	50	)and B(	39	);
	C	(	2547	)	<= A(	51	)and B(	39	);
	C	(	2548	)	<= A(	52	)and B(	39	);
	C	(	2549	)	<= A(	53	)and B(	39	);
	C	(	2550	)	<= A(	54	)and B(	39	);
	C	(	2551	)	<= A(	55	)and B(	39	);
	C	(	2552	)	<= A(	56	)and B(	39	);
	C	(	2553	)	<= A(	57	)and B(	39	);
	C	(	2554	)	<= A(	58	)and B(	39	);
	C	(	2555	)	<= A(	59	)and B(	39	);
	C	(	2556	)	<= A(	60	)and B(	39	);
	C	(	2557	)	<= A(	61	)and B(	39	);
	C	(	2558	)	<= A(	62	)and B(	39	);
	C	(	2559	)	<= A(	63	)and B(	39	);

	C	(	2560	)	<= A(	0	)and B(	40	);
	C	(	2561	)	<= A(	1	)and B(	40	);
	C	(	2562	)	<= A(	2	)and B(	40	);
	C	(	2563	)	<= A(	3	)and B(	40	);
	C	(	2564	)	<= A(	4	)and B(	40	);
	C	(	2565	)	<= A(	5	)and B(	40	);
	C	(	2566	)	<= A(	6	)and B(	40	);
	C	(	2567	)	<= A(	7	)and B(	40	);
	C	(	2568	)	<= A(	8	)and B(	40	);
	C	(	2569	)	<= A(	9	)and B(	40	);
	C	(	2570	)	<= A(	10	)and B(	40	);
	C	(	2571	)	<= A(	11	)and B(	40	);
	C	(	2572	)	<= A(	12	)and B(	40	);
	C	(	2573	)	<= A(	13	)and B(	40	);
	C	(	2574	)	<= A(	14	)and B(	40	);
	C	(	2575	)	<= A(	15	)and B(	40	);
	C	(	2576	)	<= A(	16	)and B(	40	);
	C	(	2577	)	<= A(	17	)and B(	40	);
	C	(	2578	)	<= A(	18	)and B(	40	);
	C	(	2579	)	<= A(	19	)and B(	40	);
	C	(	2580	)	<= A(	20	)and B(	40	);
	C	(	2581	)	<= A(	21	)and B(	40	);
	C	(	2582	)	<= A(	22	)and B(	40	);
	C	(	2583	)	<= A(	23	)and B(	40	);
	C	(	2584	)	<= A(	24	)and B(	40	);
	C	(	2585	)	<= A(	25	)and B(	40	);
	C	(	2586	)	<= A(	26	)and B(	40	);
	C	(	2587	)	<= A(	27	)and B(	40	);
	C	(	2588	)	<= A(	28	)and B(	40	);
	C	(	2589	)	<= A(	29	)and B(	40	);
	C	(	2590	)	<= A(	30	)and B(	40	);
	C	(	2591	)	<= A(	31	)and B(	40	);
	C	(	2592	)	<= A(	32	)and B(	40	);
	C	(	2593	)	<= A(	33	)and B(	40	);
	C	(	2594	)	<= A(	34	)and B(	40	);
	C	(	2595	)	<= A(	35	)and B(	40	);
	C	(	2596	)	<= A(	36	)and B(	40	);
	C	(	2597	)	<= A(	37	)and B(	40	);
	C	(	2598	)	<= A(	38	)and B(	40	);
	C	(	2599	)	<= A(	39	)and B(	40	);
	C	(	2600	)	<= A(	40	)and B(	40	);
	C	(	2601	)	<= A(	41	)and B(	40	);
	C	(	2602	)	<= A(	42	)and B(	40	);
	C	(	2603	)	<= A(	43	)and B(	40	);
	C	(	2604	)	<= A(	44	)and B(	40	);
	C	(	2605	)	<= A(	45	)and B(	40	);
	C	(	2606	)	<= A(	46	)and B(	40	);
	C	(	2607	)	<= A(	47	)and B(	40	);
	C	(	2608	)	<= A(	48	)and B(	40	);
	C	(	2609	)	<= A(	49	)and B(	40	);
	C	(	2610	)	<= A(	50	)and B(	40	);
	C	(	2611	)	<= A(	51	)and B(	40	);
	C	(	2612	)	<= A(	52	)and B(	40	);
	C	(	2613	)	<= A(	53	)and B(	40	);
	C	(	2614	)	<= A(	54	)and B(	40	);
	C	(	2615	)	<= A(	55	)and B(	40	);
	C	(	2616	)	<= A(	56	)and B(	40	);
	C	(	2617	)	<= A(	57	)and B(	40	);
	C	(	2618	)	<= A(	58	)and B(	40	);
	C	(	2619	)	<= A(	59	)and B(	40	);
	C	(	2620	)	<= A(	60	)and B(	40	);
	C	(	2621	)	<= A(	61	)and B(	40	);
	C	(	2622	)	<= A(	62	)and B(	40	);
	C	(	2623	)	<= A(	63	)and B(	40	);

	C	(	2624	)	<= A(	0	)and B(	41	);
	C	(	2625	)	<= A(	1	)and B(	41	);
	C	(	2626	)	<= A(	2	)and B(	41	);
	C	(	2627	)	<= A(	3	)and B(	41	);
	C	(	2628	)	<= A(	4	)and B(	41	);
	C	(	2629	)	<= A(	5	)and B(	41	);
	C	(	2630	)	<= A(	6	)and B(	41	);
	C	(	2631	)	<= A(	7	)and B(	41	);
	C	(	2632	)	<= A(	8	)and B(	41	);
	C	(	2633	)	<= A(	9	)and B(	41	);
	C	(	2634	)	<= A(	10	)and B(	41	);
	C	(	2635	)	<= A(	11	)and B(	41	);
	C	(	2636	)	<= A(	12	)and B(	41	);
	C	(	2637	)	<= A(	13	)and B(	41	);
	C	(	2638	)	<= A(	14	)and B(	41	);
	C	(	2639	)	<= A(	15	)and B(	41	);
	C	(	2640	)	<= A(	16	)and B(	41	);
	C	(	2641	)	<= A(	17	)and B(	41	);
	C	(	2642	)	<= A(	18	)and B(	41	);
	C	(	2643	)	<= A(	19	)and B(	41	);
	C	(	2644	)	<= A(	20	)and B(	41	);
	C	(	2645	)	<= A(	21	)and B(	41	);
	C	(	2646	)	<= A(	22	)and B(	41	);
	C	(	2647	)	<= A(	23	)and B(	41	);
	C	(	2648	)	<= A(	24	)and B(	41	);
	C	(	2649	)	<= A(	25	)and B(	41	);
	C	(	2650	)	<= A(	26	)and B(	41	);
	C	(	2651	)	<= A(	27	)and B(	41	);
	C	(	2652	)	<= A(	28	)and B(	41	);
	C	(	2653	)	<= A(	29	)and B(	41	);
	C	(	2654	)	<= A(	30	)and B(	41	);
	C	(	2655	)	<= A(	31	)and B(	41	);
	C	(	2656	)	<= A(	32	)and B(	41	);
	C	(	2657	)	<= A(	33	)and B(	41	);
	C	(	2658	)	<= A(	34	)and B(	41	);
	C	(	2659	)	<= A(	35	)and B(	41	);
	C	(	2660	)	<= A(	36	)and B(	41	);
	C	(	2661	)	<= A(	37	)and B(	41	);
	C	(	2662	)	<= A(	38	)and B(	41	);
	C	(	2663	)	<= A(	39	)and B(	41	);
	C	(	2664	)	<= A(	40	)and B(	41	);
	C	(	2665	)	<= A(	41	)and B(	41	);
	C	(	2666	)	<= A(	42	)and B(	41	);
	C	(	2667	)	<= A(	43	)and B(	41	);
	C	(	2668	)	<= A(	44	)and B(	41	);
	C	(	2669	)	<= A(	45	)and B(	41	);
	C	(	2670	)	<= A(	46	)and B(	41	);
	C	(	2671	)	<= A(	47	)and B(	41	);
	C	(	2672	)	<= A(	48	)and B(	41	);
	C	(	2673	)	<= A(	49	)and B(	41	);
	C	(	2674	)	<= A(	50	)and B(	41	);
	C	(	2675	)	<= A(	51	)and B(	41	);
	C	(	2676	)	<= A(	52	)and B(	41	);
	C	(	2677	)	<= A(	53	)and B(	41	);
	C	(	2678	)	<= A(	54	)and B(	41	);
	C	(	2679	)	<= A(	55	)and B(	41	);
	C	(	2680	)	<= A(	56	)and B(	41	);
	C	(	2681	)	<= A(	57	)and B(	41	);
	C	(	2682	)	<= A(	58	)and B(	41	);
	C	(	2683	)	<= A(	59	)and B(	41	);
	C	(	2684	)	<= A(	60	)and B(	41	);
	C	(	2685	)	<= A(	61	)and B(	41	);
	C	(	2686	)	<= A(	62	)and B(	41	);
	C	(	2687	)	<= A(	63	)and B(	41	);

	C	(	2688	)	<= A(	0	)and B(	42	);
	C	(	2689	)	<= A(	1	)and B(	42	);
	C	(	2690	)	<= A(	2	)and B(	42	);
	C	(	2691	)	<= A(	3	)and B(	42	);
	C	(	2692	)	<= A(	4	)and B(	42	);
	C	(	2693	)	<= A(	5	)and B(	42	);
	C	(	2694	)	<= A(	6	)and B(	42	);
	C	(	2695	)	<= A(	7	)and B(	42	);
	C	(	2696	)	<= A(	8	)and B(	42	);
	C	(	2697	)	<= A(	9	)and B(	42	);
	C	(	2698	)	<= A(	10	)and B(	42	);
	C	(	2699	)	<= A(	11	)and B(	42	);
	C	(	2700	)	<= A(	12	)and B(	42	);
	C	(	2701	)	<= A(	13	)and B(	42	);
	C	(	2702	)	<= A(	14	)and B(	42	);
	C	(	2703	)	<= A(	15	)and B(	42	);
	C	(	2704	)	<= A(	16	)and B(	42	);
	C	(	2705	)	<= A(	17	)and B(	42	);
	C	(	2706	)	<= A(	18	)and B(	42	);
	C	(	2707	)	<= A(	19	)and B(	42	);
	C	(	2708	)	<= A(	20	)and B(	42	);
	C	(	2709	)	<= A(	21	)and B(	42	);
	C	(	2710	)	<= A(	22	)and B(	42	);
	C	(	2711	)	<= A(	23	)and B(	42	);
	C	(	2712	)	<= A(	24	)and B(	42	);
	C	(	2713	)	<= A(	25	)and B(	42	);
	C	(	2714	)	<= A(	26	)and B(	42	);
	C	(	2715	)	<= A(	27	)and B(	42	);
	C	(	2716	)	<= A(	28	)and B(	42	);
	C	(	2717	)	<= A(	29	)and B(	42	);
	C	(	2718	)	<= A(	30	)and B(	42	);
	C	(	2719	)	<= A(	31	)and B(	42	);
	C	(	2720	)	<= A(	32	)and B(	42	);
	C	(	2721	)	<= A(	33	)and B(	42	);
	C	(	2722	)	<= A(	34	)and B(	42	);
	C	(	2723	)	<= A(	35	)and B(	42	);
	C	(	2724	)	<= A(	36	)and B(	42	);
	C	(	2725	)	<= A(	37	)and B(	42	);
	C	(	2726	)	<= A(	38	)and B(	42	);
	C	(	2727	)	<= A(	39	)and B(	42	);
	C	(	2728	)	<= A(	40	)and B(	42	);
	C	(	2729	)	<= A(	41	)and B(	42	);
	C	(	2730	)	<= A(	42	)and B(	42	);
	C	(	2731	)	<= A(	43	)and B(	42	);
	C	(	2732	)	<= A(	44	)and B(	42	);
	C	(	2733	)	<= A(	45	)and B(	42	);
	C	(	2734	)	<= A(	46	)and B(	42	);
	C	(	2735	)	<= A(	47	)and B(	42	);
	C	(	2736	)	<= A(	48	)and B(	42	);
	C	(	2737	)	<= A(	49	)and B(	42	);
	C	(	2738	)	<= A(	50	)and B(	42	);
	C	(	2739	)	<= A(	51	)and B(	42	);
	C	(	2740	)	<= A(	52	)and B(	42	);
	C	(	2741	)	<= A(	53	)and B(	42	);
	C	(	2742	)	<= A(	54	)and B(	42	);
	C	(	2743	)	<= A(	55	)and B(	42	);
	C	(	2744	)	<= A(	56	)and B(	42	);
	C	(	2745	)	<= A(	57	)and B(	42	);
	C	(	2746	)	<= A(	58	)and B(	42	);
	C	(	2747	)	<= A(	59	)and B(	42	);
	C	(	2748	)	<= A(	60	)and B(	42	);
	C	(	2749	)	<= A(	61	)and B(	42	);
	C	(	2750	)	<= A(	62	)and B(	42	);
	C	(	2751	)	<= A(	63	)and B(	42	);

 	C	(	2752	)	<= A(	0	)and B(	43	);
	C	(	2753	)	<= A(	1	)and B(	43	);
	C	(	2754	)	<= A(	2	)and B(	43	);
	C	(	2755	)	<= A(	3	)and B(	43	);
	C	(	2756	)	<= A(	4	)and B(	43	);
	C	(	2757	)	<= A(	5	)and B(	43	);
	C	(	2758	)	<= A(	6	)and B(	43	);
	C	(	2759	)	<= A(	7	)and B(	43	);
	C	(	2760	)	<= A(	8	)and B(	43	);
	C	(	2761	)	<= A(	9	)and B(	43	);
	C	(	2762	)	<= A(	10	)and B(	43	);
	C	(	2763	)	<= A(	11	)and B(	43	);
	C	(	2764	)	<= A(	12	)and B(	43	);
	C	(	2765	)	<= A(	13	)and B(	43	);
	C	(	2766	)	<= A(	14	)and B(	43	);
	C	(	2767	)	<= A(	15	)and B(	43	);
	C	(	2768	)	<= A(	16	)and B(	43	);
	C	(	2769	)	<= A(	17	)and B(	43	);
	C	(	2770	)	<= A(	18	)and B(	43	);
	C	(	2771	)	<= A(	19	)and B(	43	);
	C	(	2772	)	<= A(	20	)and B(	43	);
	C	(	2773	)	<= A(	21	)and B(	43	);
	C	(	2774	)	<= A(	22	)and B(	43	);
	C	(	2775	)	<= A(	23	)and B(	43	);
	C	(	2776	)	<= A(	24	)and B(	43	);
	C	(	2777	)	<= A(	25	)and B(	43	);
	C	(	2778	)	<= A(	26	)and B(	43	);
	C	(	2779	)	<= A(	27	)and B(	43	);
	C	(	2780	)	<= A(	28	)and B(	43	);
	C	(	2781	)	<= A(	29	)and B(	43	);
	C	(	2782	)	<= A(	30	)and B(	43	);
	C	(	2783	)	<= A(	31	)and B(	43	);
	C	(	2784	)	<= A(	32	)and B(	43	);
	C	(	2785	)	<= A(	33	)and B(	43	);
	C	(	2786	)	<= A(	34	)and B(	43	);
	C	(	2787	)	<= A(	35	)and B(	43	);
	C	(	2788	)	<= A(	36	)and B(	43	);
	C	(	2789	)	<= A(	37	)and B(	43	);
	C	(	2790	)	<= A(	38	)and B(	43	);
	C	(	2791	)	<= A(	39	)and B(	43	);
	C	(	2792	)	<= A(	40	)and B(	43	);
	C	(	2793	)	<= A(	41	)and B(	43	);
	C	(	2794	)	<= A(	42	)and B(	43	);
	C	(	2795	)	<= A(	43	)and B(	43	);
	C	(	2796	)	<= A(	44	)and B(	43	);
	C	(	2797	)	<= A(	45	)and B(	43	);
	C	(	2798	)	<= A(	46	)and B(	43	);
	C	(	2799	)	<= A(	47	)and B(	43	);
	C	(	2800	)	<= A(	48	)and B(	43	);
	C	(	2801	)	<= A(	49	)and B(	43	);
	C	(	2802	)	<= A(	50	)and B(	43	);
	C	(	2803	)	<= A(	51	)and B(	43	);
	C	(	2804	)	<= A(	52	)and B(	43	);
	C	(	2805	)	<= A(	53	)and B(	43	);
	C	(	2806	)	<= A(	54	)and B(	43	);
	C	(	2807	)	<= A(	55	)and B(	43	);
	C	(	2808	)	<= A(	56	)and B(	43	);
	C	(	2809	)	<= A(	57	)and B(	43	);
	C	(	2810	)	<= A(	58	)and B(	43	);
	C	(	2811	)	<= A(	59	)and B(	43	);
	C	(	2812	)	<= A(	60	)and B(	43	);
	C	(	2813	)	<= A(	61	)and B(	43	);
	C	(	2814	)	<= A(	62	)and B(	43	);
	C	(	2815	)	<= A(	63	)and B(	43	);

	C	(	2816	)	<= A(	0	)and B(	44	);
	C	(	2817	)	<= A(	1	)and B(	44	);
	C	(	2818	)	<= A(	2	)and B(	44	);
	C	(	2819	)	<= A(	3	)and B(	44	);
	C	(	2820	)	<= A(	4	)and B(	44	);
	C	(	2821	)	<= A(	5	)and B(	44	);
	C	(	2822	)	<= A(	6	)and B(	44	);
	C	(	2823	)	<= A(	7	)and B(	44	);
	C	(	2824	)	<= A(	8	)and B(	44	);
	C	(	2825	)	<= A(	9	)and B(	44	);
	C	(	2826	)	<= A(	10	)and B(	44	);
	C	(	2827	)	<= A(	11	)and B(	44	);
	C	(	2828	)	<= A(	12	)and B(	44	);
	C	(	2829	)	<= A(	13	)and B(	44	);
	C	(	2830	)	<= A(	14	)and B(	44	);
	C	(	2831	)	<= A(	15	)and B(	44	);
	C	(	2832	)	<= A(	16	)and B(	44	);
	C	(	2833	)	<= A(	17	)and B(	44	);
	C	(	2834	)	<= A(	18	)and B(	44	);
	C	(	2835	)	<= A(	19	)and B(	44	);
	C	(	2836	)	<= A(	20	)and B(	44	);
	C	(	2837	)	<= A(	21	)and B(	44	);
	C	(	2838	)	<= A(	22	)and B(	44	);
	C	(	2839	)	<= A(	23	)and B(	44	);
	C	(	2840	)	<= A(	24	)and B(	44	);
	C	(	2841	)	<= A(	25	)and B(	44	);
	C	(	2842	)	<= A(	26	)and B(	44	);
	C	(	2843	)	<= A(	27	)and B(	44	);
	C	(	2844	)	<= A(	28	)and B(	44	);
	C	(	2845	)	<= A(	29	)and B(	44	);
	C	(	2846	)	<= A(	30	)and B(	44	);
	C	(	2847	)	<= A(	31	)and B(	44	);
	C	(	2848	)	<= A(	32	)and B(	44	);
	C	(	2849	)	<= A(	33	)and B(	44	);
	C	(	2850	)	<= A(	34	)and B(	44	);
	C	(	2851	)	<= A(	35	)and B(	44	);
	C	(	2852	)	<= A(	36	)and B(	44	);
	C	(	2853	)	<= A(	37	)and B(	44	);
	C	(	2854	)	<= A(	38	)and B(	44	);
	C	(	2855	)	<= A(	39	)and B(	44	);
	C	(	2856	)	<= A(	40	)and B(	44	);
	C	(	2857	)	<= A(	41	)and B(	44	);
	C	(	2858	)	<= A(	42	)and B(	44	);
	C	(	2859	)	<= A(	43	)and B(	44	);
	C	(	2860	)	<= A(	44	)and B(	44	);
	C	(	2861	)	<= A(	45	)and B(	44	);
	C	(	2862	)	<= A(	46	)and B(	44	);
	C	(	2863	)	<= A(	47	)and B(	44	);
	C	(	2864	)	<= A(	48	)and B(	44	);
	C	(	2865	)	<= A(	49	)and B(	44	);
	C	(	2866	)	<= A(	50	)and B(	44	);
	C	(	2867	)	<= A(	51	)and B(	44	);
	C	(	2868	)	<= A(	52	)and B(	44	);
	C	(	2869	)	<= A(	53	)and B(	44	);
	C	(	2870	)	<= A(	54	)and B(	44	);
	C	(	2871	)	<= A(	55	)and B(	44	);
	C	(	2872	)	<= A(	56	)and B(	44	);
	C	(	2873	)	<= A(	57	)and B(	44	);
	C	(	2874	)	<= A(	58	)and B(	44	);
	C	(	2875	)	<= A(	59	)and B(	44	);
	C	(	2876	)	<= A(	60	)and B(	44	);
	C	(	2877	)	<= A(	61	)and B(	44	);
	C	(	2878	)	<= A(	62	)and B(	44	);
	C	(	2879	)	<= A(	63	)and B(	44	);

	C	(	2880	)	<= A(	0	)and B(	45	);
	C	(	2881	)	<= A(	1	)and B(	45	);
	C	(	2882	)	<= A(	2	)and B(	45	);
	C	(	2883	)	<= A(	3	)and B(	45	);
	C	(	2884	)	<= A(	4	)and B(	45	);
	C	(	2885	)	<= A(	5	)and B(	45	);
	C	(	2886	)	<= A(	6	)and B(	45	);
	C	(	2887	)	<= A(	7	)and B(	45	);
	C	(	2888	)	<= A(	8	)and B(	45	);
	C	(	2889	)	<= A(	9	)and B(	45	);
	C	(	2890	)	<= A(	10	)and B(	45	);
	C	(	2891	)	<= A(	11	)and B(	45	);
	C	(	2892	)	<= A(	12	)and B(	45	);
	C	(	2893	)	<= A(	13	)and B(	45	);
	C	(	2894	)	<= A(	14	)and B(	45	);
	C	(	2895	)	<= A(	15	)and B(	45	);
	C	(	2896	)	<= A(	16	)and B(	45	);
	C	(	2897	)	<= A(	17	)and B(	45	);
	C	(	2898	)	<= A(	18	)and B(	45	);
	C	(	2899	)	<= A(	19	)and B(	45	);
	C	(	2900	)	<= A(	20	)and B(	45	);
	C	(	2901	)	<= A(	21	)and B(	45	);
	C	(	2902	)	<= A(	22	)and B(	45	);
	C	(	2903	)	<= A(	23	)and B(	45	);
	C	(	2904	)	<= A(	24	)and B(	45	);
	C	(	2905	)	<= A(	25	)and B(	45	);
	C	(	2906	)	<= A(	26	)and B(	45	);
	C	(	2907	)	<= A(	27	)and B(	45	);
	C	(	2908	)	<= A(	28	)and B(	45	);
	C	(	2909	)	<= A(	29	)and B(	45	);
	C	(	2910	)	<= A(	30	)and B(	45	);
	C	(	2911	)	<= A(	31	)and B(	45	);
	C	(	2912	)	<= A(	32	)and B(	45	);
	C	(	2913	)	<= A(	33	)and B(	45	);
	C	(	2914	)	<= A(	34	)and B(	45	);
	C	(	2915	)	<= A(	35	)and B(	45	);
	C	(	2916	)	<= A(	36	)and B(	45	);
	C	(	2917	)	<= A(	37	)and B(	45	);
	C	(	2918	)	<= A(	38	)and B(	45	);
	C	(	2919	)	<= A(	39	)and B(	45	);
	C	(	2920	)	<= A(	40	)and B(	45	);
	C	(	2921	)	<= A(	41	)and B(	45	);
	C	(	2922	)	<= A(	42	)and B(	45	);
	C	(	2923	)	<= A(	43	)and B(	45	);
	C	(	2924	)	<= A(	44	)and B(	45	);
	C	(	2925	)	<= A(	45	)and B(	45	);
	C	(	2926	)	<= A(	46	)and B(	45	);
	C	(	2927	)	<= A(	47	)and B(	45	);
	C	(	2928	)	<= A(	48	)and B(	45	);
	C	(	2929	)	<= A(	49	)and B(	45	);
	C	(	2930	)	<= A(	50	)and B(	45	);
	C	(	2931	)	<= A(	51	)and B(	45	);
	C	(	2932	)	<= A(	52	)and B(	45	);
	C	(	2933	)	<= A(	53	)and B(	45	);
	C	(	2934	)	<= A(	54	)and B(	45	);
	C	(	2935	)	<= A(	55	)and B(	45	);
	C	(	2936	)	<= A(	56	)and B(	45	);
	C	(	2937	)	<= A(	57	)and B(	45	);
	C	(	2938	)	<= A(	58	)and B(	45	);
	C	(	2939	)	<= A(	59	)and B(	45	);
	C	(	2940	)	<= A(	60	)and B(	45	);
	C	(	2941	)	<= A(	61	)and B(	45	);
	C	(	2942	)	<= A(	62	)and B(	45	);
	C	(	2943	)	<= A(	63	)and B(	45	);


	C	(	2944	)	<= A(	0	)and B(	46	);
	C	(	2945	)	<= A(	1	)and B(	46	);
	C	(	2946	)	<= A(	2	)and B(	46	);
	C	(	2947	)	<= A(	3	)and B(	46	);
	C	(	2948	)	<= A(	4	)and B(	46	);
	C	(	2949	)	<= A(	5	)and B(	46	);
	C	(	2950	)	<= A(	6	)and B(	46	);
	C	(	2951	)	<= A(	7	)and B(	46	);
	C	(	2952	)	<= A(	8	)and B(	46	);
	C	(	2953	)	<= A(	9	)and B(	46	);
	C	(	2954	)	<= A(	10	)and B(	46	);
	C	(	2955	)	<= A(	11	)and B(	46	);
	C	(	2956	)	<= A(	12	)and B(	46	);
	C	(	2957	)	<= A(	13	)and B(	46	);
	C	(	2958	)	<= A(	14	)and B(	46	);
	C	(	2959	)	<= A(	15	)and B(	46	);
	C	(	2960	)	<= A(	16	)and B(	46	);
	C	(	2961	)	<= A(	17	)and B(	46	);
	C	(	2962	)	<= A(	18	)and B(	46	);
	C	(	2963	)	<= A(	19	)and B(	46	);
	C	(	2964	)	<= A(	20	)and B(	46	);
	C	(	2965	)	<= A(	21	)and B(	46	);
	C	(	2966	)	<= A(	22	)and B(	46	);
	C	(	2967	)	<= A(	23	)and B(	46	);
	C	(	2968	)	<= A(	24	)and B(	46	);
	C	(	2969	)	<= A(	25	)and B(	46	);
	C	(	2970	)	<= A(	26	)and B(	46	);
	C	(	2971	)	<= A(	27	)and B(	46	);
	C	(	2972	)	<= A(	28	)and B(	46	);
	C	(	2973	)	<= A(	29	)and B(	46	);
	C	(	2974	)	<= A(	30	)and B(	46	);
	C	(	2975	)	<= A(	31	)and B(	46	);
	C	(	2976	)	<= A(	32	)and B(	46	);
	C	(	2977	)	<= A(	33	)and B(	46	);
	C	(	2978	)	<= A(	34	)and B(	46	);
	C	(	2979	)	<= A(	35	)and B(	46	);
	C	(	2980	)	<= A(	36	)and B(	46	);
	C	(	2981	)	<= A(	37	)and B(	46	);
	C	(	2982	)	<= A(	38	)and B(	46	);
	C	(	2983	)	<= A(	39	)and B(	46	);
	C	(	2984	)	<= A(	40	)and B(	46	);
	C	(	2985	)	<= A(	41	)and B(	46	);
	C	(	2986	)	<= A(	42	)and B(	46	);
	C	(	2987	)	<= A(	43	)and B(	46	);
	C	(	2988	)	<= A(	44	)and B(	46	);
	C	(	2989	)	<= A(	45	)and B(	46	);
	C	(	2990	)	<= A(	46	)and B(	46	);
	C	(	2991	)	<= A(	47	)and B(	46	);
	C	(	2992	)	<= A(	48	)and B(	46	);
	C	(	2993	)	<= A(	49	)and B(	46	);
	C	(	2994	)	<= A(	50	)and B(	46	);
	C	(	2995	)	<= A(	51	)and B(	46	);
	C	(	2996	)	<= A(	52	)and B(	46	);
	C	(	2997	)	<= A(	53	)and B(	46	);
	C	(	2998	)	<= A(	54	)and B(	46	);
	C	(	2999	)	<= A(	55	)and B(	46	);
	C	(	3000	)	<= A(	56	)and B(	46	);
	C	(	3001	)	<= A(	57	)and B(	46	);
	C	(	3002	)	<= A(	58	)and B(	46	);
	C	(	3003	)	<= A(	59	)and B(	46	);
	C	(	3004	)	<= A(	60	)and B(	46	);
	C	(	3005	)	<= A(	61	)and B(	46	);
	C	(	3006	)	<= A(	62	)and B(	46	);
	C	(	3007	)	<= A(	63	)and B(	46	);

	C	(	3008	)	<= A(	0	)and B(	47	);
	C	(	3009	)	<= A(	1	)and B(	47	);
	C	(	3010	)	<= A(	2	)and B(	47	);
	C	(	3011	)	<= A(	3	)and B(	47	);
	C	(	3012	)	<= A(	4	)and B(	47	);
	C	(	3013	)	<= A(	5	)and B(	47	);
	C	(	3014	)	<= A(	6	)and B(	47	);
	C	(	3015	)	<= A(	7	)and B(	47	);
	C	(	3016	)	<= A(	8	)and B(	47	);
	C	(	3017	)	<= A(	9	)and B(	47	);
	C	(	3018	)	<= A(	10	)and B(	47	);
	C	(	3019	)	<= A(	11	)and B(	47	);
	C	(	3020	)	<= A(	12	)and B(	47	);
	C	(	3021	)	<= A(	13	)and B(	47	);
	C	(	3022	)	<= A(	14	)and B(	47	);
	C	(	3023	)	<= A(	15	)and B(	47	);
	C	(	3024	)	<= A(	16	)and B(	47	);
	C	(	3025	)	<= A(	17	)and B(	47	);
	C	(	3026	)	<= A(	18	)and B(	47	);
	C	(	3027	)	<= A(	19	)and B(	47	);
	C	(	3028	)	<= A(	20	)and B(	47	);
	C	(	3029	)	<= A(	21	)and B(	47	);
	C	(	3030	)	<= A(	22	)and B(	47	);
	C	(	3031	)	<= A(	23	)and B(	47	);
	C	(	3032	)	<= A(	24	)and B(	47	);
	C	(	3033	)	<= A(	25	)and B(	47	);
	C	(	3034	)	<= A(	26	)and B(	47	);
	C	(	3035	)	<= A(	27	)and B(	47	);
	C	(	3036	)	<= A(	28	)and B(	47	);
	C	(	3037	)	<= A(	29	)and B(	47	);
	C	(	3038	)	<= A(	30	)and B(	47	);
	C	(	3039	)	<= A(	31	)and B(	47	);
	C	(	3040	)	<= A(	32	)and B(	47	);
	C	(	3041	)	<= A(	33	)and B(	47	);
	C	(	3042	)	<= A(	34	)and B(	47	);
	C	(	3043	)	<= A(	35	)and B(	47	);
	C	(	3044	)	<= A(	36	)and B(	47	);
	C	(	3045	)	<= A(	37	)and B(	47	);
	C	(	3046	)	<= A(	38	)and B(	47	);
	C	(	3047	)	<= A(	39	)and B(	47	);
	C	(	3048	)	<= A(	40	)and B(	47	);
	C	(	3049	)	<= A(	41	)and B(	47	);
	C	(	3050	)	<= A(	42	)and B(	47	);
	C	(	3051	)	<= A(	43	)and B(	47	);
	C	(	3052	)	<= A(	44	)and B(	47	);
	C	(	3053	)	<= A(	45	)and B(	47	);
	C	(	3054	)	<= A(	46	)and B(	47	);
	C	(	3055	)	<= A(	47	)and B(	47	);
	C	(	3056	)	<= A(	48	)and B(	47	);
	C	(	3057	)	<= A(	49	)and B(	47	);
	C	(	3058	)	<= A(	50	)and B(	47	);
	C	(	3059	)	<= A(	51	)and B(	47	);
	C	(	3060	)	<= A(	52	)and B(	47	);
	C	(	3061	)	<= A(	53	)and B(	47	);
	C	(	3062	)	<= A(	54	)and B(	47	);
	C	(	3063	)	<= A(	55	)and B(	47	);
	C	(	3064	)	<= A(	56	)and B(	47	);
	C	(	3065	)	<= A(	57	)and B(	47	);
	C	(	3066	)	<= A(	58	)and B(	47	);
	C	(	3067	)	<= A(	59	)and B(	47	);
	C	(	3068	)	<= A(	60	)and B(	47	);
	C	(	3069	)	<= A(	61	)and B(	47	);
	C	(	3070	)	<= A(	62	)and B(	47	);
	C	(	3071	)	<= A(	63	)and B(	47	);

	C	(	3072	)	<= A(	0	)and B(	48	);
	C	(	3073	)	<= A(	1	)and B(	48	);
	C	(	3074	)	<= A(	2	)and B(	48	);
	C	(	3075	)	<= A(	3	)and B(	48	);
	C	(	3076	)	<= A(	4	)and B(	48	);
	C	(	3077	)	<= A(	5	)and B(	48	);
	C	(	3078	)	<= A(	6	)and B(	48	);
	C	(	3079	)	<= A(	7	)and B(	48	);
	C	(	3080	)	<= A(	8	)and B(	48	);
	C	(	3081	)	<= A(	9	)and B(	48	);
	C	(	3082	)	<= A(	10	)and B(	48	);
	C	(	3083	)	<= A(	11	)and B(	48	);
	C	(	3084	)	<= A(	12	)and B(	48	);
	C	(	3085	)	<= A(	13	)and B(	48	);
	C	(	3086	)	<= A(	14	)and B(	48	);
	C	(	3087	)	<= A(	15	)and B(	48	);
	C	(	3088	)	<= A(	16	)and B(	48	);
	C	(	3089	)	<= A(	17	)and B(	48	);
	C	(	3090	)	<= A(	18	)and B(	48	);
	C	(	3091	)	<= A(	19	)and B(	48	);
	C	(	3092	)	<= A(	20	)and B(	48	);
	C	(	3093	)	<= A(	21	)and B(	48	);
	C	(	3094	)	<= A(	22	)and B(	48	);
	C	(	3095	)	<= A(	23	)and B(	48	);
	C	(	3096	)	<= A(	24	)and B(	48	);
	C	(	3097	)	<= A(	25	)and B(	48	);
	C	(	3098	)	<= A(	26	)and B(	48	);
	C	(	3099	)	<= A(	27	)and B(	48	);
	C	(	3100	)	<= A(	28	)and B(	48	);
	C	(	3101	)	<= A(	29	)and B(	48	);
	C	(	3102	)	<= A(	30	)and B(	48	);
	C	(	3103	)	<= A(	31	)and B(	48	);
	C	(	3104	)	<= A(	32	)and B(	48	);
	C	(	3105	)	<= A(	33	)and B(	48	);
	C	(	3106	)	<= A(	34	)and B(	48	);
	C	(	3107	)	<= A(	35	)and B(	48	);
	C	(	3108	)	<= A(	36	)and B(	48	);
	C	(	3109	)	<= A(	37	)and B(	48	);
	C	(	3110	)	<= A(	38	)and B(	48	);
	C	(	3111	)	<= A(	39	)and B(	48	);
	C	(	3112	)	<= A(	40	)and B(	48	);
	C	(	3113	)	<= A(	41	)and B(	48	);
	C	(	3114	)	<= A(	42	)and B(	48	);
	C	(	3115	)	<= A(	43	)and B(	48	);
	C	(	3116	)	<= A(	44	)and B(	48	);
	C	(	3117	)	<= A(	45	)and B(	48	);
	C	(	3118	)	<= A(	46	)and B(	48	);
	C	(	3119	)	<= A(	47	)and B(	48	);
	C	(	3120	)	<= A(	48	)and B(	48	);
	C	(	3121	)	<= A(	49	)and B(	48	);
	C	(	3122	)	<= A(	50	)and B(	48	);
	C	(	3123	)	<= A(	51	)and B(	48	);
	C	(	3124	)	<= A(	52	)and B(	48	);
	C	(	3125	)	<= A(	53	)and B(	48	);
	C	(	3126	)	<= A(	54	)and B(	48	);
	C	(	3127	)	<= A(	55	)and B(	48	);
	C	(	3128	)	<= A(	56	)and B(	48	);
	C	(	3129	)	<= A(	57	)and B(	48	);
	C	(	3130	)	<= A(	58	)and B(	48	);
	C	(	3131	)	<= A(	59	)and B(	48	);
	C	(	3132	)	<= A(	60	)and B(	48	);
	C	(	3133	)	<= A(	61	)and B(	48	);
	C	(	3134	)	<= A(	62	)and B(	48	);
	C	(	3135	)	<= A(	63	)and B(	48	);

	C	(	3136	)	<= A(	0	)and B(	49	);
	C	(	3137	)	<= A(	1	)and B(	49	);
	C	(	3138	)	<= A(	2	)and B(	49	);
	C	(	3139	)	<= A(	3	)and B(	49	);
	C	(	3140	)	<= A(	4	)and B(	49	);
	C	(	3141	)	<= A(	5	)and B(	49	);
	C	(	3142	)	<= A(	6	)and B(	49	);
	C	(	3143	)	<= A(	7	)and B(	49	);
	C	(	3144	)	<= A(	8	)and B(	49	);
	C	(	3145	)	<= A(	9	)and B(	49	);
	C	(	3146	)	<= A(	10	)and B(	49	);
	C	(	3147	)	<= A(	11	)and B(	49	);
	C	(	3148	)	<= A(	12	)and B(	49	);
	C	(	3149	)	<= A(	13	)and B(	49	);
	C	(	3150	)	<= A(	14	)and B(	49	);
	C	(	3151	)	<= A(	15	)and B(	49	);
	C	(	3152	)	<= A(	16	)and B(	49	);
	C	(	3153	)	<= A(	17	)and B(	49	);
	C	(	3154	)	<= A(	18	)and B(	49	);
	C	(	3155	)	<= A(	19	)and B(	49	);
	C	(	3156	)	<= A(	20	)and B(	49	);
	C	(	3157	)	<= A(	21	)and B(	49	);
	C	(	3158	)	<= A(	22	)and B(	49	);
	C	(	3159	)	<= A(	23	)and B(	49	);
	C	(	3160	)	<= A(	24	)and B(	49	);
	C	(	3161	)	<= A(	25	)and B(	49	);
	C	(	3162	)	<= A(	26	)and B(	49	);
	C	(	3163	)	<= A(	27	)and B(	49	);
	C	(	3164	)	<= A(	28	)and B(	49	);
	C	(	3165	)	<= A(	29	)and B(	49	);
	C	(	3166	)	<= A(	30	)and B(	49	);
	C	(	3167	)	<= A(	31	)and B(	49	);
	C	(	3168	)	<= A(	32	)and B(	49	);
	C	(	3169	)	<= A(	33	)and B(	49	);
	C	(	3170	)	<= A(	34	)and B(	49	);
	C	(	3171	)	<= A(	35	)and B(	49	);
	C	(	3172	)	<= A(	36	)and B(	49	);
	C	(	3173	)	<= A(	37	)and B(	49	);
	C	(	3174	)	<= A(	38	)and B(	49	);
	C	(	3175	)	<= A(	39	)and B(	49	);
	C	(	3176	)	<= A(	40	)and B(	49	);
	C	(	3177	)	<= A(	41	)and B(	49	);
	C	(	3178	)	<= A(	42	)and B(	49	);
	C	(	3179	)	<= A(	43	)and B(	49	);
	C	(	3180	)	<= A(	44	)and B(	49	);
	C	(	3181	)	<= A(	45	)and B(	49	);
	C	(	3182	)	<= A(	46	)and B(	49	);
	C	(	3183	)	<= A(	47	)and B(	49	);
	C	(	3184	)	<= A(	48	)and B(	49	);
	C	(	3185	)	<= A(	49	)and B(	49	);
	C	(	3186	)	<= A(	50	)and B(	49	);
	C	(	3187	)	<= A(	51	)and B(	49	);
	C	(	3188	)	<= A(	52	)and B(	49	);
	C	(	3189	)	<= A(	53	)and B(	49	);
	C	(	3190	)	<= A(	54	)and B(	49	);
	C	(	3191	)	<= A(	55	)and B(	49	);
	C	(	3192	)	<= A(	56	)and B(	49	);
	C	(	3193	)	<= A(	57	)and B(	49	);
	C	(	3194	)	<= A(	58	)and B(	49	);
	C	(	3195	)	<= A(	59	)and B(	49	);
	C	(	3196	)	<= A(	60	)and B(	49	);
	C	(	3197	)	<= A(	61	)and B(	49	);
	C	(	3198	)	<= A(	62	)and B(	49	);
	C	(	3199	)	<= A(	63	)and B(	49	);


	C	(	3200	)	<= A(	0	)and B(	50	);
	C	(	3201	)	<= A(	1	)and B(	50	);
	C	(	3202	)	<= A(	2	)and B(	50	);
	C	(	3203	)	<= A(	3	)and B(	50	);
	C	(	3204	)	<= A(	4	)and B(	50	);
	C	(	3205	)	<= A(	5	)and B(	50	);
	C	(	3206	)	<= A(	6	)and B(	50	);
	C	(	3207	)	<= A(	7	)and B(	50	);
	C	(	3208	)	<= A(	8	)and B(	50	);
	C	(	3209	)	<= A(	9	)and B(	50	);
	C	(	3210	)	<= A(	10	)and B(	50	);
	C	(	3211	)	<= A(	11	)and B(	50	);
	C	(	3212	)	<= A(	12	)and B(	50	);
	C	(	3213	)	<= A(	13	)and B(	50	);
	C	(	3214	)	<= A(	14	)and B(	50	);
	C	(	3215	)	<= A(	15	)and B(	50	);
	C	(	3216	)	<= A(	16	)and B(	50	);
	C	(	3217	)	<= A(	17	)and B(	50	);
	C	(	3218	)	<= A(	18	)and B(	50	);
	C	(	3219	)	<= A(	19	)and B(	50	);
	C	(	3220	)	<= A(	20	)and B(	50	);
	C	(	3221	)	<= A(	21	)and B(	50	);
	C	(	3222	)	<= A(	22	)and B(	50	);
	C	(	3223	)	<= A(	23	)and B(	50	);
	C	(	3224	)	<= A(	24	)and B(	50	);
	C	(	3225	)	<= A(	25	)and B(	50	);
	C	(	3226	)	<= A(	26	)and B(	50	);
	C	(	3227	)	<= A(	27	)and B(	50	);
	C	(	3228	)	<= A(	28	)and B(	50	);
	C	(	3229	)	<= A(	29	)and B(	50	);
	C	(	3230	)	<= A(	30	)and B(	50	);
	C	(	3231	)	<= A(	31	)and B(	50	);
	C	(	3232	)	<= A(	32	)and B(	50	);
	C	(	3233	)	<= A(	33	)and B(	50	);
	C	(	3234	)	<= A(	34	)and B(	50	);
	C	(	3235	)	<= A(	35	)and B(	50	);
	C	(	3236	)	<= A(	36	)and B(	50	);
	C	(	3237	)	<= A(	37	)and B(	50	);
	C	(	3238	)	<= A(	38	)and B(	50	);
	C	(	3239	)	<= A(	39	)and B(	50	);
	C	(	3240	)	<= A(	40	)and B(	50	);
	C	(	3241	)	<= A(	41	)and B(	50	);
	C	(	3242	)	<= A(	42	)and B(	50	);
	C	(	3243	)	<= A(	43	)and B(	50	);
	C	(	3244	)	<= A(	44	)and B(	50	);
	C	(	3245	)	<= A(	45	)and B(	50	);
	C	(	3246	)	<= A(	46	)and B(	50	);
	C	(	3247	)	<= A(	47	)and B(	50	);
	C	(	3248	)	<= A(	48	)and B(	50	);
	C	(	3249	)	<= A(	49	)and B(	50	);
	C	(	3250	)	<= A(	50	)and B(	50	);
	C	(	3251	)	<= A(	51	)and B(	50	);
	C	(	3252	)	<= A(	52	)and B(	50	);
	C	(	3253	)	<= A(	53	)and B(	50	);
	C	(	3254	)	<= A(	54	)and B(	50	);
	C	(	3255	)	<= A(	55	)and B(	50	);
	C	(	3256	)	<= A(	56	)and B(	50	);
	C	(	3257	)	<= A(	57	)and B(	50	);
	C	(	3258	)	<= A(	58	)and B(	50	);
	C	(	3259	)	<= A(	59	)and B(	50	);
	C	(	3260	)	<= A(	60	)and B(	50	);
	C	(	3261	)	<= A(	61	)and B(	50	);
	C	(	3262	)	<= A(	62	)and B(	50	);
	C	(	3263	)	<= A(	63	)and B(	50	);

	C	(	3264	)	<= A(	0	)and B(	51	);
	C	(	3265	)	<= A(	1	)and B(	51	);
	C	(	3266	)	<= A(	2	)and B(	51	);
	C	(	3267	)	<= A(	3	)and B(	51	);
	C	(	3268	)	<= A(	4	)and B(	51	);
	C	(	3269	)	<= A(	5	)and B(	51	);
	C	(	3270	)	<= A(	6	)and B(	51	);
	C	(	3271	)	<= A(	7	)and B(	51	);
	C	(	3272	)	<= A(	8	)and B(	51	);
	C	(	3273	)	<= A(	9	)and B(	51	);
	C	(	3274	)	<= A(	10	)and B(	51	);
	C	(	3275	)	<= A(	11	)and B(	51	);
	C	(	3276	)	<= A(	12	)and B(	51	);
	C	(	3277	)	<= A(	13	)and B(	51	);
	C	(	3278	)	<= A(	14	)and B(	51	);
	C	(	3279	)	<= A(	15	)and B(	51	);
	C	(	3280	)	<= A(	16	)and B(	51	);
	C	(	3281	)	<= A(	17	)and B(	51	);
	C	(	3282	)	<= A(	18	)and B(	51	);
	C	(	3283	)	<= A(	19	)and B(	51	);
	C	(	3284	)	<= A(	20	)and B(	51	);
	C	(	3285	)	<= A(	21	)and B(	51	);
	C	(	3286	)	<= A(	22	)and B(	51	);
	C	(	3287	)	<= A(	23	)and B(	51	);
	C	(	3288	)	<= A(	24	)and B(	51	);
	C	(	3289	)	<= A(	25	)and B(	51	);
	C	(	3290	)	<= A(	26	)and B(	51	);
	C	(	3291	)	<= A(	27	)and B(	51	);
	C	(	3292	)	<= A(	28	)and B(	51	);
	C	(	3293	)	<= A(	29	)and B(	51	);
	C	(	3294	)	<= A(	30	)and B(	51	);
	C	(	3295	)	<= A(	31	)and B(	51	);
	C	(	3296	)	<= A(	32	)and B(	51	);
	C	(	3297	)	<= A(	33	)and B(	51	);
	C	(	3298	)	<= A(	34	)and B(	51	);
	C	(	3299	)	<= A(	35	)and B(	51	);
	C	(	3300	)	<= A(	36	)and B(	51	);
	C	(	3301	)	<= A(	37	)and B(	51	);
	C	(	3302	)	<= A(	38	)and B(	51	);
	C	(	3303	)	<= A(	39	)and B(	51	);
	C	(	3304	)	<= A(	40	)and B(	51	);
	C	(	3305	)	<= A(	41	)and B(	51	);
	C	(	3306	)	<= A(	42	)and B(	51	);
	C	(	3307	)	<= A(	43	)and B(	51	);
	C	(	3308	)	<= A(	44	)and B(	51	);
	C	(	3309	)	<= A(	45	)and B(	51	);
	C	(	3310	)	<= A(	46	)and B(	51	);
	C	(	3311	)	<= A(	47	)and B(	51	);
	C	(	3312	)	<= A(	48	)and B(	51	);
	C	(	3313	)	<= A(	49	)and B(	51	);
	C	(	3314	)	<= A(	50	)and B(	51	);
	C	(	3315	)	<= A(	51	)and B(	51	);
	C	(	3316	)	<= A(	52	)and B(	51	);
	C	(	3317	)	<= A(	53	)and B(	51	);
	C	(	3318	)	<= A(	54	)and B(	51	);
	C	(	3319	)	<= A(	55	)and B(	51	);
	C	(	3320	)	<= A(	56	)and B(	51	);
	C	(	3321	)	<= A(	57	)and B(	51	);
	C	(	3322	)	<= A(	58	)and B(	51	);
	C	(	3323	)	<= A(	59	)and B(	51	);
	C	(	3324	)	<= A(	60	)and B(	51	);
	C	(	3325	)	<= A(	61	)and B(	51	);
	C	(	3326	)	<= A(	62	)and B(	51	);
	C	(	3327	)	<= A(	63	)and B(	51	);

	C	(	3328	)	<= A(	0	)and B(	52	);
	C	(	3329	)	<= A(	1	)and B(	52	);
	C	(	3330	)	<= A(	2	)and B(	52	);
	C	(	3331	)	<= A(	3	)and B(	52	);
	C	(	3332	)	<= A(	4	)and B(	52	);
	C	(	3333	)	<= A(	5	)and B(	52	);
	C	(	3334	)	<= A(	6	)and B(	52	);
	C	(	3335	)	<= A(	7	)and B(	52	);
	C	(	3336	)	<= A(	8	)and B(	52	);
	C	(	3337	)	<= A(	9	)and B(	52	);
	C	(	3338	)	<= A(	10	)and B(	52	);
	C	(	3339	)	<= A(	11	)and B(	52	);
	C	(	3340	)	<= A(	12	)and B(	52	);
	C	(	3341	)	<= A(	13	)and B(	52	);
	C	(	3342	)	<= A(	14	)and B(	52	);
	C	(	3343	)	<= A(	15	)and B(	52	);
	C	(	3344	)	<= A(	16	)and B(	52	);
	C	(	3345	)	<= A(	17	)and B(	52	);
	C	(	3346	)	<= A(	18	)and B(	52	);
	C	(	3347	)	<= A(	19	)and B(	52	);
	C	(	3348	)	<= A(	20	)and B(	52	);
	C	(	3349	)	<= A(	21	)and B(	52	);
	C	(	3350	)	<= A(	22	)and B(	52	);
	C	(	3351	)	<= A(	23	)and B(	52	);
	C	(	3352	)	<= A(	24	)and B(	52	);
	C	(	3353	)	<= A(	25	)and B(	52	);
	C	(	3354	)	<= A(	26	)and B(	52	);
	C	(	3355	)	<= A(	27	)and B(	52	);
	C	(	3356	)	<= A(	28	)and B(	52	);
	C	(	3357	)	<= A(	29	)and B(	52	);
	C	(	3358	)	<= A(	30	)and B(	52	);
	C	(	3359	)	<= A(	31	)and B(	52	);
	C	(	3360	)	<= A(	32	)and B(	52	);
	C	(	3361	)	<= A(	33	)and B(	52	);
	C	(	3362	)	<= A(	34	)and B(	52	);
	C	(	3363	)	<= A(	35	)and B(	52	);
	C	(	3364	)	<= A(	36	)and B(	52	);
	C	(	3365	)	<= A(	37	)and B(	52	);
	C	(	3366	)	<= A(	38	)and B(	52	);
	C	(	3367	)	<= A(	39	)and B(	52	);
	C	(	3368	)	<= A(	40	)and B(	52	);
	C	(	3369	)	<= A(	41	)and B(	52	);
	C	(	3370	)	<= A(	42	)and B(	52	);
	C	(	3371	)	<= A(	43	)and B(	52	);
	C	(	3372	)	<= A(	44	)and B(	52	);
	C	(	3373	)	<= A(	45	)and B(	52	);
	C	(	3374	)	<= A(	46	)and B(	52	);
	C	(	3375	)	<= A(	47	)and B(	52	);
	C	(	3376	)	<= A(	48	)and B(	52	);
	C	(	3377	)	<= A(	49	)and B(	52	);
	C	(	3378	)	<= A(	50	)and B(	52	);
	C	(	3379	)	<= A(	51	)and B(	52	);
	C	(	3380	)	<= A(	52	)and B(	52	);
	C	(	3381	)	<= A(	53	)and B(	52	);
	C	(	3382	)	<= A(	54	)and B(	52	);
	C	(	3383	)	<= A(	55	)and B(	52	);
	C	(	3384	)	<= A(	56	)and B(	52	);
	C	(	3385	)	<= A(	57	)and B(	52	);
	C	(	3386	)	<= A(	58	)and B(	52	);
	C	(	3387	)	<= A(	59	)and B(	52	);
	C	(	3388	)	<= A(	60	)and B(	52	);
	C	(	3389	)	<= A(	61	)and B(	52	);
	C	(	3390	)	<= A(	62	)and B(	52	);
	C	(	3391	)	<= A(	63	)and B(	52	);

	C	(	3392	)	<= A(	0	)and B(	53	);
	C	(	3393	)	<= A(	1	)and B(	53	);
	C	(	3394	)	<= A(	2	)and B(	53	);
	C	(	3395	)	<= A(	3	)and B(	53	);
	C	(	3396	)	<= A(	4	)and B(	53	);
	C	(	3397	)	<= A(	5	)and B(	53	);
	C	(	3398	)	<= A(	6	)and B(	53	);
	C	(	3399	)	<= A(	7	)and B(	53	);
	C	(	3400	)	<= A(	8	)and B(	53	);
	C	(	3401	)	<= A(	9	)and B(	53	);
	C	(	3402	)	<= A(	10	)and B(	53	);
	C	(	3403	)	<= A(	11	)and B(	53	);
	C	(	3404	)	<= A(	12	)and B(	53	);
	C	(	3405	)	<= A(	13	)and B(	53	);
	C	(	3406	)	<= A(	14	)and B(	53	);
	C	(	3407	)	<= A(	15	)and B(	53	);
	C	(	3408	)	<= A(	16	)and B(	53	);
	C	(	3409	)	<= A(	17	)and B(	53	);
	C	(	3410	)	<= A(	18	)and B(	53	);
	C	(	3411	)	<= A(	19	)and B(	53	);
	C	(	3412	)	<= A(	20	)and B(	53	);
	C	(	3413	)	<= A(	21	)and B(	53	);
	C	(	3414	)	<= A(	22	)and B(	53	);
	C	(	3415	)	<= A(	23	)and B(	53	);
	C	(	3416	)	<= A(	24	)and B(	53	);
	C	(	3417	)	<= A(	25	)and B(	53	);
	C	(	3418	)	<= A(	26	)and B(	53	);
	C	(	3419	)	<= A(	27	)and B(	53	);
	C	(	3420	)	<= A(	28	)and B(	53	);
	C	(	3421	)	<= A(	29	)and B(	53	);
	C	(	3422	)	<= A(	30	)and B(	53	);
	C	(	3423	)	<= A(	31	)and B(	53	);
	C	(	3424	)	<= A(	32	)and B(	53	);
	C	(	3425	)	<= A(	33	)and B(	53	);
	C	(	3426	)	<= A(	34	)and B(	53	);
	C	(	3427	)	<= A(	35	)and B(	53	);
	C	(	3428	)	<= A(	36	)and B(	53	);
	C	(	3429	)	<= A(	37	)and B(	53	);
	C	(	3430	)	<= A(	38	)and B(	53	);
	C	(	3431	)	<= A(	39	)and B(	53	);
	C	(	3432	)	<= A(	40	)and B(	53	);
	C	(	3433	)	<= A(	41	)and B(	53	);
	C	(	3434	)	<= A(	42	)and B(	53	);
	C	(	3435	)	<= A(	43	)and B(	53	);
	C	(	3436	)	<= A(	44	)and B(	53	);
	C	(	3437	)	<= A(	45	)and B(	53	);
	C	(	3438	)	<= A(	46	)and B(	53	);
	C	(	3439	)	<= A(	47	)and B(	53	);
	C	(	3440	)	<= A(	48	)and B(	53	);
	C	(	3441	)	<= A(	49	)and B(	53	);
	C	(	3442	)	<= A(	50	)and B(	53	);
	C	(	3443	)	<= A(	51	)and B(	53	);
	C	(	3444	)	<= A(	52	)and B(	53	);
	C	(	3445	)	<= A(	53	)and B(	53	);
	C	(	3446	)	<= A(	54	)and B(	53	);
	C	(	3447	)	<= A(	55	)and B(	53	);
	C	(	3448	)	<= A(	56	)and B(	53	);
	C	(	3449	)	<= A(	57	)and B(	53	);
	C	(	3450	)	<= A(	58	)and B(	53	);
	C	(	3451	)	<= A(	59	)and B(	53	);
	C	(	3452	)	<= A(	60	)and B(	53	);
	C	(	3453	)	<= A(	61	)and B(	53	);
	C	(	3454	)	<= A(	62	)and B(	53	);
	C	(	3455	)	<= A(	63	)and B(	53	);

	C	(	3456	)	<= A(	0	)and B(	54	);
	C	(	3457	)	<= A(	1	)and B(	54	);
	C	(	3458	)	<= A(	2	)and B(	54	);
	C	(	3459	)	<= A(	3	)and B(	54	);
	C	(	3460	)	<= A(	4	)and B(	54	);
	C	(	3461	)	<= A(	5	)and B(	54	);
	C	(	3462	)	<= A(	6	)and B(	54	);
	C	(	3463	)	<= A(	7	)and B(	54	);
	C	(	3464	)	<= A(	8	)and B(	54	);
	C	(	3465	)	<= A(	9	)and B(	54	);
	C	(	3466	)	<= A(	10	)and B(	54	);
	C	(	3467	)	<= A(	11	)and B(	54	);
	C	(	3468	)	<= A(	12	)and B(	54	);
	C	(	3469	)	<= A(	13	)and B(	54	);
	C	(	3470	)	<= A(	14	)and B(	54	);
	C	(	3471	)	<= A(	15	)and B(	54	);
	C	(	3472	)	<= A(	16	)and B(	54	);
	C	(	3473	)	<= A(	17	)and B(	54	);
	C	(	3474	)	<= A(	18	)and B(	54	);
	C	(	3475	)	<= A(	19	)and B(	54	);
	C	(	3476	)	<= A(	20	)and B(	54	);
	C	(	3477	)	<= A(	21	)and B(	54	);
	C	(	3478	)	<= A(	22	)and B(	54	);
	C	(	3479	)	<= A(	23	)and B(	54	);
	C	(	3480	)	<= A(	24	)and B(	54	);
	C	(	3481	)	<= A(	25	)and B(	54	);
	C	(	3482	)	<= A(	26	)and B(	54	);
	C	(	3483	)	<= A(	27	)and B(	54	);
	C	(	3484	)	<= A(	28	)and B(	54	);
	C	(	3485	)	<= A(	29	)and B(	54	);
	C	(	3486	)	<= A(	30	)and B(	54	);
	C	(	3487	)	<= A(	31	)and B(	54	);
	C	(	3488	)	<= A(	32	)and B(	54	);
	C	(	3489	)	<= A(	33	)and B(	54	);
	C	(	3490	)	<= A(	34	)and B(	54	);
	C	(	3491	)	<= A(	35	)and B(	54	);
	C	(	3492	)	<= A(	36	)and B(	54	);
	C	(	3493	)	<= A(	37	)and B(	54	);
	C	(	3494	)	<= A(	38	)and B(	54	);
	C	(	3495	)	<= A(	39	)and B(	54	);
	C	(	3496	)	<= A(	40	)and B(	54	);
	C	(	3497	)	<= A(	41	)and B(	54	);
	C	(	3498	)	<= A(	42	)and B(	54	);
	C	(	3499	)	<= A(	43	)and B(	54	);
	C	(	3500	)	<= A(	44	)and B(	54	);
	C	(	3501	)	<= A(	45	)and B(	54	);
	C	(	3502	)	<= A(	46	)and B(	54	);
	C	(	3503	)	<= A(	47	)and B(	54	);
	C	(	3504	)	<= A(	48	)and B(	54	);
	C	(	3505	)	<= A(	49	)and B(	54	);
	C	(	3506	)	<= A(	50	)and B(	54	);
	C	(	3507	)	<= A(	51	)and B(	54	);
	C	(	3508	)	<= A(	52	)and B(	54	);
	C	(	3509	)	<= A(	53	)and B(	54	);
	C	(	3510	)	<= A(	54	)and B(	54	);
	C	(	3511	)	<= A(	55	)and B(	54	);
	C	(	3512	)	<= A(	56	)and B(	54	);
	C	(	3513	)	<= A(	57	)and B(	54	);
	C	(	3514	)	<= A(	58	)and B(	54	);
	C	(	3515	)	<= A(	59	)and B(	54	);
	C	(	3516	)	<= A(	60	)and B(	54	);
	C	(	3517	)	<= A(	61	)and B(	54	);
	C	(	3518	)	<= A(	62	)and B(	54	);
	C	(	3519	)	<= A(	63	)and B(	54	);

	C	(	3520	)	<= A(	0	)and B(	55	);
	C	(	3521	)	<= A(	1	)and B(	55	);
	C	(	3522	)	<= A(	2	)and B(	55	);
	C	(	3523	)	<= A(	3	)and B(	55	);
	C	(	3524	)	<= A(	4	)and B(	55	);
	C	(	3525	)	<= A(	5	)and B(	55	);
	C	(	3526	)	<= A(	6	)and B(	55	);
	C	(	3527	)	<= A(	7	)and B(	55	);
	C	(	3528	)	<= A(	8	)and B(	55	);
	C	(	3529	)	<= A(	9	)and B(	55	);
	C	(	3530	)	<= A(	10	)and B(	55	);
	C	(	3531	)	<= A(	11	)and B(	55	);
	C	(	3532	)	<= A(	12	)and B(	55	);
	C	(	3533	)	<= A(	13	)and B(	55	);
	C	(	3534	)	<= A(	14	)and B(	55	);
	C	(	3535	)	<= A(	15	)and B(	55	);
	C	(	3536	)	<= A(	16	)and B(	55	);
	C	(	3537	)	<= A(	17	)and B(	55	);
	C	(	3538	)	<= A(	18	)and B(	55	);
	C	(	3539	)	<= A(	19	)and B(	55	);
	C	(	3540	)	<= A(	20	)and B(	55	);
	C	(	3541	)	<= A(	21	)and B(	55	);
	C	(	3542	)	<= A(	22	)and B(	55	);
	C	(	3543	)	<= A(	23	)and B(	55	);
	C	(	3544	)	<= A(	24	)and B(	55	);
	C	(	3545	)	<= A(	25	)and B(	55	);
	C	(	3546	)	<= A(	26	)and B(	55	);
	C	(	3547	)	<= A(	27	)and B(	55	);
	C	(	3548	)	<= A(	28	)and B(	55	);
	C	(	3549	)	<= A(	29	)and B(	55	);
	C	(	3550	)	<= A(	30	)and B(	55	);
	C	(	3551	)	<= A(	31	)and B(	55	);
	C	(	3552	)	<= A(	32	)and B(	55	);
	C	(	3553	)	<= A(	33	)and B(	55	);
	C	(	3554	)	<= A(	34	)and B(	55	);
	C	(	3555	)	<= A(	35	)and B(	55	);
	C	(	3556	)	<= A(	36	)and B(	55	);
	C	(	3557	)	<= A(	37	)and B(	55	);
	C	(	3558	)	<= A(	38	)and B(	55	);
	C	(	3559	)	<= A(	39	)and B(	55	);
	C	(	3560	)	<= A(	40	)and B(	55	);
	C	(	3561	)	<= A(	41	)and B(	55	);
	C	(	3562	)	<= A(	42	)and B(	55	);
	C	(	3563	)	<= A(	43	)and B(	55	);
	C	(	3564	)	<= A(	44	)and B(	55	);
	C	(	3565	)	<= A(	45	)and B(	55	);
	C	(	3566	)	<= A(	46	)and B(	55	);
	C	(	3567	)	<= A(	47	)and B(	55	);
	C	(	3568	)	<= A(	48	)and B(	55	);
	C	(	3569	)	<= A(	49	)and B(	55	);
	C	(	3570	)	<= A(	50	)and B(	55	);
	C	(	3571	)	<= A(	51	)and B(	55	);
	C	(	3572	)	<= A(	52	)and B(	55	);
	C	(	3573	)	<= A(	53	)and B(	55	);
	C	(	3574	)	<= A(	54	)and B(	55	);
	C	(	3575	)	<= A(	55	)and B(	55	);
	C	(	3576	)	<= A(	56	)and B(	55	);
	C	(	3577	)	<= A(	57	)and B(	55	);
	C	(	3578	)	<= A(	58	)and B(	55	);
	C	(	3579	)	<= A(	59	)and B(	55	);
	C	(	3580	)	<= A(	60	)and B(	55	);
	C	(	3581	)	<= A(	61	)and B(	55	);
	C	(	3582	)	<= A(	62	)and B(	55	);
	C	(	3583	)	<= A(	63	)and B(	55	);

	C	(	3584	)	<= A(	0	)and B(	56	);
	C	(	3585	)	<= A(	1	)and B(	56	);
	C	(	3586	)	<= A(	2	)and B(	56	);
	C	(	3587	)	<= A(	3	)and B(	56	);
	C	(	3588	)	<= A(	4	)and B(	56	);
	C	(	3589	)	<= A(	5	)and B(	56	);
	C	(	3590	)	<= A(	6	)and B(	56	);
	C	(	3591	)	<= A(	7	)and B(	56	);
	C	(	3592	)	<= A(	8	)and B(	56	);
	C	(	3593	)	<= A(	9	)and B(	56	);
	C	(	3594	)	<= A(	10	)and B(	56	);
	C	(	3595	)	<= A(	11	)and B(	56	);
	C	(	3596	)	<= A(	12	)and B(	56	);
	C	(	3597	)	<= A(	13	)and B(	56	);
	C	(	3598	)	<= A(	14	)and B(	56	);
	C	(	3599	)	<= A(	15	)and B(	56	);
	C	(	3600	)	<= A(	16	)and B(	56	);
	C	(	3601	)	<= A(	17	)and B(	56	);
	C	(	3602	)	<= A(	18	)and B(	56	);
	C	(	3603	)	<= A(	19	)and B(	56	);
	C	(	3604	)	<= A(	20	)and B(	56	);
	C	(	3605	)	<= A(	21	)and B(	56	);
	C	(	3606	)	<= A(	22	)and B(	56	);
	C	(	3607	)	<= A(	23	)and B(	56	);
	C	(	3608	)	<= A(	24	)and B(	56	);
	C	(	3609	)	<= A(	25	)and B(	56	);
	C	(	3610	)	<= A(	26	)and B(	56	);
	C	(	3611	)	<= A(	27	)and B(	56	);
	C	(	3612	)	<= A(	28	)and B(	56	);
	C	(	3613	)	<= A(	29	)and B(	56	);
	C	(	3614	)	<= A(	30	)and B(	56	);
	C	(	3615	)	<= A(	31	)and B(	56	);
	C	(	3616	)	<= A(	32	)and B(	56	);
	C	(	3617	)	<= A(	33	)and B(	56	);
	C	(	3618	)	<= A(	34	)and B(	56	);
	C	(	3619	)	<= A(	35	)and B(	56	);
	C	(	3620	)	<= A(	36	)and B(	56	);
	C	(	3621	)	<= A(	37	)and B(	56	);
	C	(	3622	)	<= A(	38	)and B(	56	);
	C	(	3623	)	<= A(	39	)and B(	56	);
	C	(	3624	)	<= A(	40	)and B(	56	);
	C	(	3625	)	<= A(	41	)and B(	56	);
	C	(	3626	)	<= A(	42	)and B(	56	);
	C	(	3627	)	<= A(	43	)and B(	56	);
	C	(	3628	)	<= A(	44	)and B(	56	);
	C	(	3629	)	<= A(	45	)and B(	56	);
	C	(	3630	)	<= A(	46	)and B(	56	);
	C	(	3631	)	<= A(	47	)and B(	56	);
	C	(	3632	)	<= A(	48	)and B(	56	);
	C	(	3633	)	<= A(	49	)and B(	56	);
	C	(	3634	)	<= A(	50	)and B(	56	);
	C	(	3635	)	<= A(	51	)and B(	56	);
	C	(	3636	)	<= A(	52	)and B(	56	);
	C	(	3637	)	<= A(	53	)and B(	56	);
	C	(	3638	)	<= A(	54	)and B(	56	);
	C	(	3639	)	<= A(	55	)and B(	56	);
	C	(	3640	)	<= A(	56	)and B(	56	);
	C	(	3641	)	<= A(	57	)and B(	56	);
	C	(	3642	)	<= A(	58	)and B(	56	);
	C	(	3643	)	<= A(	59	)and B(	56	);
	C	(	3644	)	<= A(	60	)and B(	56	);
	C	(	3645	)	<= A(	61	)and B(	56	);
	C	(	3646	)	<= A(	62	)and B(	56	);
	C	(	3647	)	<= A(	63	)and B(	56	);

	C	(	3648	)	<= A(	0	)and B(	57	);
	C	(	3649	)	<= A(	1	)and B(	57	);
	C	(	3650	)	<= A(	2	)and B(	57	);
	C	(	3651	)	<= A(	3	)and B(	57	);
	C	(	3652	)	<= A(	4	)and B(	57	);
	C	(	3653	)	<= A(	5	)and B(	57	);
	C	(	3654	)	<= A(	6	)and B(	57	);
	C	(	3655	)	<= A(	7	)and B(	57	);
	C	(	3656	)	<= A(	8	)and B(	57	);
	C	(	3657	)	<= A(	9	)and B(	57	);
	C	(	3658	)	<= A(	10	)and B(	57	);
	C	(	3659	)	<= A(	11	)and B(	57	);
	C	(	3660	)	<= A(	12	)and B(	57	);
	C	(	3661	)	<= A(	13	)and B(	57	);
	C	(	3662	)	<= A(	14	)and B(	57	);
	C	(	3663	)	<= A(	15	)and B(	57	);
	C	(	3664	)	<= A(	16	)and B(	57	);
	C	(	3665	)	<= A(	17	)and B(	57	);
	C	(	3666	)	<= A(	18	)and B(	57	);
	C	(	3667	)	<= A(	19	)and B(	57	);
	C	(	3668	)	<= A(	20	)and B(	57	);
	C	(	3669	)	<= A(	21	)and B(	57	);
	C	(	3670	)	<= A(	22	)and B(	57	);
	C	(	3671	)	<= A(	23	)and B(	57	);
	C	(	3672	)	<= A(	24	)and B(	57	);
	C	(	3673	)	<= A(	25	)and B(	57	);
	C	(	3674	)	<= A(	26	)and B(	57	);
	C	(	3675	)	<= A(	27	)and B(	57	);
	C	(	3676	)	<= A(	28	)and B(	57	);
	C	(	3677	)	<= A(	29	)and B(	57	);
	C	(	3678	)	<= A(	30	)and B(	57	);
	C	(	3679	)	<= A(	31	)and B(	57	);
	C	(	3680	)	<= A(	32	)and B(	57	);
	C	(	3681	)	<= A(	33	)and B(	57	);
	C	(	3682	)	<= A(	34	)and B(	57	);
	C	(	3683	)	<= A(	35	)and B(	57	);
	C	(	3684	)	<= A(	36	)and B(	57	);
	C	(	3685	)	<= A(	37	)and B(	57	);
	C	(	3686	)	<= A(	38	)and B(	57	);
	C	(	3687	)	<= A(	39	)and B(	57	);
	C	(	3688	)	<= A(	40	)and B(	57	);
	C	(	3689	)	<= A(	41	)and B(	57	);
	C	(	3690	)	<= A(	42	)and B(	57	);
	C	(	3691	)	<= A(	43	)and B(	57	);
	C	(	3692	)	<= A(	44	)and B(	57	);
	C	(	3693	)	<= A(	45	)and B(	57	);
	C	(	3694	)	<= A(	46	)and B(	57	);
	C	(	3695	)	<= A(	47	)and B(	57	);
	C	(	3696	)	<= A(	48	)and B(	57	);
	C	(	3697	)	<= A(	49	)and B(	57	);
	C	(	3698	)	<= A(	50	)and B(	57	);
	C	(	3699	)	<= A(	51	)and B(	57	);
	C	(	3700	)	<= A(	52	)and B(	57	);
	C	(	3701	)	<= A(	53	)and B(	57	);
	C	(	3702	)	<= A(	54	)and B(	57	);
	C	(	3703	)	<= A(	55	)and B(	57	);
	C	(	3704	)	<= A(	56	)and B(	57	);
	C	(	3705	)	<= A(	57	)and B(	57	);
	C	(	3706	)	<= A(	58	)and B(	57	);
	C	(	3707	)	<= A(	59	)and B(	57	);
	C	(	3708	)	<= A(	60	)and B(	57	);
	C	(	3709	)	<= A(	61	)and B(	57	);
	C	(	3710	)	<= A(	62	)and B(	57	);
	C	(	3711	)	<= A(	63	)and B(	57	);

	C	(	3712	)	<= A(	0	)and B(	58	);
	C	(	3713	)	<= A(	1	)and B(	58	);
	C	(	3714	)	<= A(	2	)and B(	58	);
	C	(	3715	)	<= A(	3	)and B(	58	);
	C	(	3716	)	<= A(	4	)and B(	58	);
	C	(	3717	)	<= A(	5	)and B(	58	);
	C	(	3718	)	<= A(	6	)and B(	58	);
	C	(	3719	)	<= A(	7	)and B(	58	);
	C	(	3720	)	<= A(	8	)and B(	58	);
	C	(	3721	)	<= A(	9	)and B(	58	);
	C	(	3722	)	<= A(	10	)and B(	58	);
	C	(	3723	)	<= A(	11	)and B(	58	);
	C	(	3724	)	<= A(	12	)and B(	58	);
	C	(	3725	)	<= A(	13	)and B(	58	);
	C	(	3726	)	<= A(	14	)and B(	58	);
	C	(	3727	)	<= A(	15	)and B(	58	);
	C	(	3728	)	<= A(	16	)and B(	58	);
	C	(	3729	)	<= A(	17	)and B(	58	);
	C	(	3730	)	<= A(	18	)and B(	58	);
	C	(	3731	)	<= A(	19	)and B(	58	);
	C	(	3732	)	<= A(	20	)and B(	58	);
	C	(	3733	)	<= A(	21	)and B(	58	);
	C	(	3734	)	<= A(	22	)and B(	58	);
	C	(	3735	)	<= A(	23	)and B(	58	);
	C	(	3736	)	<= A(	24	)and B(	58	);
	C	(	3737	)	<= A(	25	)and B(	58	);
	C	(	3738	)	<= A(	26	)and B(	58	);
	C	(	3739	)	<= A(	27	)and B(	58	);
	C	(	3740	)	<= A(	28	)and B(	58	);
	C	(	3741	)	<= A(	29	)and B(	58	);
	C	(	3742	)	<= A(	30	)and B(	58	);
	C	(	3743	)	<= A(	31	)and B(	58	);
	C	(	3744	)	<= A(	32	)and B(	58	);
	C	(	3745	)	<= A(	33	)and B(	58	);
	C	(	3746	)	<= A(	34	)and B(	58	);
	C	(	3747	)	<= A(	35	)and B(	58	);
	C	(	3748	)	<= A(	36	)and B(	58	);
	C	(	3749	)	<= A(	37	)and B(	58	);
	C	(	3750	)	<= A(	38	)and B(	58	);
	C	(	3751	)	<= A(	39	)and B(	58	);
	C	(	3752	)	<= A(	40	)and B(	58	);
	C	(	3753	)	<= A(	41	)and B(	58	);
	C	(	3754	)	<= A(	42	)and B(	58	);
	C	(	3755	)	<= A(	43	)and B(	58	);
	C	(	3756	)	<= A(	44	)and B(	58	);
	C	(	3757	)	<= A(	45	)and B(	58	);
	C	(	3758	)	<= A(	46	)and B(	58	);
	C	(	3759	)	<= A(	47	)and B(	58	);
	C	(	3760	)	<= A(	48	)and B(	58	);
	C	(	3761	)	<= A(	49	)and B(	58	);
	C	(	3762	)	<= A(	50	)and B(	58	);
	C	(	3763	)	<= A(	51	)and B(	58	);
	C	(	3764	)	<= A(	52	)and B(	58	);
	C	(	3765	)	<= A(	53	)and B(	58	);
	C	(	3766	)	<= A(	54	)and B(	58	);
	C	(	3767	)	<= A(	55	)and B(	58	);
	C	(	3768	)	<= A(	56	)and B(	58	);
	C	(	3769	)	<= A(	57	)and B(	58	);
	C	(	3770	)	<= A(	58	)and B(	58	);
	C	(	3771	)	<= A(	59	)and B(	58	);
	C	(	3772	)	<= A(	60	)and B(	58	);
	C	(	3773	)	<= A(	61	)and B(	58	);
	C	(	3774	)	<= A(	62	)and B(	58	);
	C	(	3775	)	<= A(	63	)and B(	58	);

	C	(	3776	)	<= A(	0	)and B(	59	);
	C	(	3777	)	<= A(	1	)and B(	59	);
	C	(	3778	)	<= A(	2	)and B(	59	);
	C	(	3779	)	<= A(	3	)and B(	59	);
	C	(	3780	)	<= A(	4	)and B(	59	);
	C	(	3781	)	<= A(	5	)and B(	59	);
	C	(	3782	)	<= A(	6	)and B(	59	);
	C	(	3783	)	<= A(	7	)and B(	59	);
	C	(	3784	)	<= A(	8	)and B(	59	);
	C	(	3785	)	<= A(	9	)and B(	59	);
	C	(	3786	)	<= A(	10	)and B(	59	);
	C	(	3787	)	<= A(	11	)and B(	59	);
	C	(	3788	)	<= A(	12	)and B(	59	);
	C	(	3789	)	<= A(	13	)and B(	59	);
	C	(	3790	)	<= A(	14	)and B(	59	);
	C	(	3791	)	<= A(	15	)and B(	59	);
	C	(	3792	)	<= A(	16	)and B(	59	);
	C	(	3793	)	<= A(	17	)and B(	59	);
	C	(	3794	)	<= A(	18	)and B(	59	);
	C	(	3795	)	<= A(	19	)and B(	59	);
	C	(	3796	)	<= A(	20	)and B(	59	);
	C	(	3797	)	<= A(	21	)and B(	59	);
	C	(	3798	)	<= A(	22	)and B(	59	);
	C	(	3799	)	<= A(	23	)and B(	59	);
	C	(	3800	)	<= A(	24	)and B(	59	);
	C	(	3801	)	<= A(	25	)and B(	59	);
	C	(	3802	)	<= A(	26	)and B(	59	);
	C	(	3803	)	<= A(	27	)and B(	59	);
	C	(	3804	)	<= A(	28	)and B(	59	);
	C	(	3805	)	<= A(	29	)and B(	59	);
	C	(	3806	)	<= A(	30	)and B(	59	);
	C	(	3807	)	<= A(	31	)and B(	59	);
	C	(	3808	)	<= A(	32	)and B(	59	);
	C	(	3809	)	<= A(	33	)and B(	59	);
	C	(	3810	)	<= A(	34	)and B(	59	);
	C	(	3811	)	<= A(	35	)and B(	59	);
	C	(	3812	)	<= A(	36	)and B(	59	);
	C	(	3813	)	<= A(	37	)and B(	59	);
	C	(	3814	)	<= A(	38	)and B(	59	);
	C	(	3815	)	<= A(	39	)and B(	59	);
	C	(	3816	)	<= A(	40	)and B(	59	);
	C	(	3817	)	<= A(	41	)and B(	59	);
	C	(	3818	)	<= A(	42	)and B(	59	);
	C	(	3819	)	<= A(	43	)and B(	59	);
	C	(	3820	)	<= A(	44	)and B(	59	);
	C	(	3821	)	<= A(	45	)and B(	59	);
	C	(	3822	)	<= A(	46	)and B(	59	);
	C	(	3823	)	<= A(	47	)and B(	59	);
	C	(	3824	)	<= A(	48	)and B(	59	);
	C	(	3825	)	<= A(	49	)and B(	59	);
	C	(	3826	)	<= A(	50	)and B(	59	);
	C	(	3827	)	<= A(	51	)and B(	59	);
	C	(	3828	)	<= A(	52	)and B(	59	);
	C	(	3829	)	<= A(	53	)and B(	59	);
	C	(	3830	)	<= A(	54	)and B(	59	);
	C	(	3831	)	<= A(	55	)and B(	59	);
	C	(	3832	)	<= A(	56	)and B(	59	);
	C	(	3833	)	<= A(	57	)and B(	59	);
	C	(	3834	)	<= A(	58	)and B(	59	);
	C	(	3835	)	<= A(	59	)and B(	59	);
	C	(	3836	)	<= A(	60	)and B(	59	);
	C	(	3837	)	<= A(	61	)and B(	59	);
	C	(	3838	)	<= A(	62	)and B(	59	);
	C	(	3839	)	<= A(	63	)and B(	59	);

	C	(	3840	)	<= A(	0	)and B(	60	);
	C	(	3841	)	<= A(	1	)and B(	60	);
	C	(	3842	)	<= A(	2	)and B(	60	);
	C	(	3843	)	<= A(	3	)and B(	60	);
	C	(	3844	)	<= A(	4	)and B(	60	);
	C	(	3845	)	<= A(	5	)and B(	60	);
	C	(	3846	)	<= A(	6	)and B(	60	);
	C	(	3847	)	<= A(	7	)and B(	60	);
	C	(	3848	)	<= A(	8	)and B(	60	);
	C	(	3849	)	<= A(	9	)and B(	60	);
	C	(	3850	)	<= A(	10	)and B(	60	);
	C	(	3851	)	<= A(	11	)and B(	60	);
	C	(	3852	)	<= A(	12	)and B(	60	);
	C	(	3853	)	<= A(	13	)and B(	60	);
	C	(	3854	)	<= A(	14	)and B(	60	);
	C	(	3855	)	<= A(	15	)and B(	60	);
	C	(	3856	)	<= A(	16	)and B(	60	);
	C	(	3857	)	<= A(	17	)and B(	60	);
	C	(	3858	)	<= A(	18	)and B(	60	);
	C	(	3859	)	<= A(	19	)and B(	60	);
	C	(	3860	)	<= A(	20	)and B(	60	);
	C	(	3861	)	<= A(	21	)and B(	60	);
	C	(	3862	)	<= A(	22	)and B(	60	);
	C	(	3863	)	<= A(	23	)and B(	60	);
	C	(	3864	)	<= A(	24	)and B(	60	);
	C	(	3865	)	<= A(	25	)and B(	60	);
	C	(	3866	)	<= A(	26	)and B(	60	);
	C	(	3867	)	<= A(	27	)and B(	60	);
	C	(	3868	)	<= A(	28	)and B(	60	);
	C	(	3869	)	<= A(	29	)and B(	60	);
	C	(	3870	)	<= A(	30	)and B(	60	);
	C	(	3871	)	<= A(	31	)and B(	60	);
	C	(	3872	)	<= A(	32	)and B(	60	);
	C	(	3873	)	<= A(	33	)and B(	60	);
	C	(	3874	)	<= A(	34	)and B(	60	);
	C	(	3875	)	<= A(	35	)and B(	60	);
	C	(	3876	)	<= A(	36	)and B(	60	);
	C	(	3877	)	<= A(	37	)and B(	60	);
	C	(	3878	)	<= A(	38	)and B(	60	);
	C	(	3879	)	<= A(	39	)and B(	60	);
	C	(	3880	)	<= A(	40	)and B(	60	);
	C	(	3881	)	<= A(	41	)and B(	60	);
	C	(	3882	)	<= A(	42	)and B(	60	);
	C	(	3883	)	<= A(	43	)and B(	60	);
	C	(	3884	)	<= A(	44	)and B(	60	);
	C	(	3885	)	<= A(	45	)and B(	60	);
	C	(	3886	)	<= A(	46	)and B(	60	);
	C	(	3887	)	<= A(	47	)and B(	60	);
	C	(	3888	)	<= A(	48	)and B(	60	);
	C	(	3889	)	<= A(	49	)and B(	60	);
	C	(	3890	)	<= A(	50	)and B(	60	);
	C	(	3891	)	<= A(	51	)and B(	60	);
	C	(	3892	)	<= A(	52	)and B(	60	);
	C	(	3893	)	<= A(	53	)and B(	60	);
	C	(	3894	)	<= A(	54	)and B(	60	);
	C	(	3895	)	<= A(	55	)and B(	60	);
	C	(	3896	)	<= A(	56	)and B(	60	);
	C	(	3897	)	<= A(	57	)and B(	60	);
	C	(	3898	)	<= A(	58	)and B(	60	);
	C	(	3899	)	<= A(	59	)and B(	60	);
	C	(	3900	)	<= A(	60	)and B(	60	);
	C	(	3901	)	<= A(	61	)and B(	60	);
	C	(	3902	)	<= A(	62	)and B(	60	);
	C	(	3903	)	<= A(	63	)and B(	60	);

	C	(	3904	)	<= A(	0	)and B(	61	);
	C	(	3905	)	<= A(	1	)and B(	61	);
	C	(	3906	)	<= A(	2	)and B(	61	);
	C	(	3907	)	<= A(	3	)and B(	61	);
	C	(	3908	)	<= A(	4	)and B(	61	);
	C	(	3909	)	<= A(	5	)and B(	61	);
	C	(	3910	)	<= A(	6	)and B(	61	);
	C	(	3911	)	<= A(	7	)and B(	61	);
	C	(	3912	)	<= A(	8	)and B(	61	);
	C	(	3913	)	<= A(	9	)and B(	61	);
	C	(	3914	)	<= A(	10	)and B(	61	);
	C	(	3915	)	<= A(	11	)and B(	61	);
	C	(	3916	)	<= A(	12	)and B(	61	);
	C	(	3917	)	<= A(	13	)and B(	61	);
	C	(	3918	)	<= A(	14	)and B(	61	);
	C	(	3919	)	<= A(	15	)and B(	61	);
	C	(	3920	)	<= A(	16	)and B(	61	);
	C	(	3921	)	<= A(	17	)and B(	61	);
	C	(	3922	)	<= A(	18	)and B(	61	);
	C	(	3923	)	<= A(	19	)and B(	61	);
	C	(	3924	)	<= A(	20	)and B(	61	);
	C	(	3925	)	<= A(	21	)and B(	61	);
	C	(	3926	)	<= A(	22	)and B(	61	);
	C	(	3927	)	<= A(	23	)and B(	61	);
	C	(	3928	)	<= A(	24	)and B(	61	);
	C	(	3929	)	<= A(	25	)and B(	61	);
	C	(	3930	)	<= A(	26	)and B(	61	);
	C	(	3931	)	<= A(	27	)and B(	61	);
	C	(	3932	)	<= A(	28	)and B(	61	);
	C	(	3933	)	<= A(	29	)and B(	61	);
	C	(	3934	)	<= A(	30	)and B(	61	);
	C	(	3935	)	<= A(	31	)and B(	61	);
	C	(	3936	)	<= A(	32	)and B(	61	);
	C	(	3937	)	<= A(	33	)and B(	61	);
	C	(	3938	)	<= A(	34	)and B(	61	);
	C	(	3939	)	<= A(	35	)and B(	61	);
	C	(	3940	)	<= A(	36	)and B(	61	);
	C	(	3941	)	<= A(	37	)and B(	61	);
	C	(	3942	)	<= A(	38	)and B(	61	);
	C	(	3943	)	<= A(	39	)and B(	61	);
	C	(	3944	)	<= A(	40	)and B(	61	);
	C	(	3945	)	<= A(	41	)and B(	61	);
	C	(	3946	)	<= A(	42	)and B(	61	);
	C	(	3947	)	<= A(	43	)and B(	61	);
	C	(	3948	)	<= A(	44	)and B(	61	);
	C	(	3949	)	<= A(	45	)and B(	61	);
	C	(	3950	)	<= A(	46	)and B(	61	);
	C	(	3951	)	<= A(	47	)and B(	61	);
	C	(	3952	)	<= A(	48	)and B(	61	);
	C	(	3953	)	<= A(	49	)and B(	61	);
	C	(	3954	)	<= A(	50	)and B(	61	);
	C	(	3955	)	<= A(	51	)and B(	61	);
	C	(	3956	)	<= A(	52	)and B(	61	);
	C	(	3957	)	<= A(	53	)and B(	61	);
	C	(	3958	)	<= A(	54	)and B(	61	);
	C	(	3959	)	<= A(	55	)and B(	61	);
	C	(	3960	)	<= A(	56	)and B(	61	);
	C	(	3961	)	<= A(	57	)and B(	61	);
	C	(	3962	)	<= A(	58	)and B(	61	);
	C	(	3963	)	<= A(	59	)and B(	61	);
	C	(	3964	)	<= A(	60	)and B(	61	);
	C	(	3965	)	<= A(	61	)and B(	61	);
	C	(	3966	)	<= A(	62	)and B(	61	);
	C	(	3967	)	<= A(	63	)and B(	61	);

	C	(	3968	)	<= A(	0	)and B(	62	);
	C	(	3969	)	<= A(	1	)and B(	62	);
	C	(	3970	)	<= A(	2	)and B(	62	);
	C	(	3971	)	<= A(	3	)and B(	62	);
	C	(	3972	)	<= A(	4	)and B(	62	);
	C	(	3973	)	<= A(	5	)and B(	62	);
	C	(	3974	)	<= A(	6	)and B(	62	);
	C	(	3975	)	<= A(	7	)and B(	62	);
	C	(	3976	)	<= A(	8	)and B(	62	);
	C	(	3977	)	<= A(	9	)and B(	62	);
	C	(	3978	)	<= A(	10	)and B(	62	);
	C	(	3979	)	<= A(	11	)and B(	62	);
	C	(	3980	)	<= A(	12	)and B(	62	);
	C	(	3981	)	<= A(	13	)and B(	62	);
	C	(	3982	)	<= A(	14	)and B(	62	);
	C	(	3983	)	<= A(	15	)and B(	62	);
	C	(	3984	)	<= A(	16	)and B(	62	);
	C	(	3985	)	<= A(	17	)and B(	62	);
	C	(	3986	)	<= A(	18	)and B(	62	);
	C	(	3987	)	<= A(	19	)and B(	62	);
	C	(	3988	)	<= A(	20	)and B(	62	);
	C	(	3989	)	<= A(	21	)and B(	62	);
	C	(	3990	)	<= A(	22	)and B(	62	);
	C	(	3991	)	<= A(	23	)and B(	62	);
	C	(	3992	)	<= A(	24	)and B(	62	);
	C	(	3993	)	<= A(	25	)and B(	62	);
	C	(	3994	)	<= A(	26	)and B(	62	);
	C	(	3995	)	<= A(	27	)and B(	62	);
	C	(	3996	)	<= A(	28	)and B(	62	);
	C	(	3997	)	<= A(	29	)and B(	62	);
	C	(	3998	)	<= A(	30	)and B(	62	);
	C	(	3999	)	<= A(	31	)and B(	62	);
	C	(	4000	)	<= A(	32	)and B(	62	);
	C	(	4001	)	<= A(	33	)and B(	62	);
	C	(	4002	)	<= A(	34	)and B(	62	);
	C	(	4003	)	<= A(	35	)and B(	62	);
	C	(	4004	)	<= A(	36	)and B(	62	);
	C	(	4005	)	<= A(	37	)and B(	62	);
	C	(	4006	)	<= A(	38	)and B(	62	);
	C	(	4007	)	<= A(	39	)and B(	62	);
	C	(	4008	)	<= A(	40	)and B(	62	);
	C	(	4009	)	<= A(	41	)and B(	62	);
	C	(	4010	)	<= A(	42	)and B(	62	);
	C	(	4011	)	<= A(	43	)and B(	62	);
	C	(	4012	)	<= A(	44	)and B(	62	);
	C	(	4013	)	<= A(	45	)and B(	62	);
	C	(	4014	)	<= A(	46	)and B(	62	);
	C	(	4015	)	<= A(	47	)and B(	62	);
	C	(	4016	)	<= A(	48	)and B(	62	);
	C	(	4017	)	<= A(	49	)and B(	62	);
	C	(	4018	)	<= A(	50	)and B(	62	);
	C	(	4019	)	<= A(	51	)and B(	62	);
	C	(	4020	)	<= A(	52	)and B(	62	);
	C	(	4021	)	<= A(	53	)and B(	62	);
	C	(	4022	)	<= A(	54	)and B(	62	);
	C	(	4023	)	<= A(	55	)and B(	62	);
	C	(	4024	)	<= A(	56	)and B(	62	);
	C	(	4025	)	<= A(	57	)and B(	62	);
	C	(	4026	)	<= A(	58	)and B(	62	);
	C	(	4027	)	<= A(	59	)and B(	62	);
	C	(	4028	)	<= A(	60	)and B(	62	);
	C	(	4029	)	<= A(	61	)and B(	62	);
	C	(	4030	)	<= A(	62	)and B(	62	);
	C	(	4031	)	<= A(	63	)and B(	62	);

	C	(	4032	)	<= A(	0	)and B(	63	);
	C	(	4033	)	<= A(	1	)and B(	63	);
	C	(	4034	)	<= A(	2	)and B(	63	);
	C	(	4035	)	<= A(	3	)and B(	63	);
	C	(	4036	)	<= A(	4	)and B(	63	);
	C	(	4037	)	<= A(	5	)and B(	63	);
	C	(	4038	)	<= A(	6	)and B(	63	);
	C	(	4039	)	<= A(	7	)and B(	63	);
	C	(	4040	)	<= A(	8	)and B(	63	);
	C	(	4041	)	<= A(	9	)and B(	63	);
	C	(	4042	)	<= A(	10	)and B(	63	);
	C	(	4043	)	<= A(	11	)and B(	63	);
	C	(	4044	)	<= A(	12	)and B(	63	);
	C	(	4045	)	<= A(	13	)and B(	63	);
	C	(	4046	)	<= A(	14	)and B(	63	);
	C	(	4047	)	<= A(	15	)and B(	63	);
	C	(	4048	)	<= A(	16	)and B(	63	);
	C	(	4049	)	<= A(	17	)and B(	63	);
	C	(	4050	)	<= A(	18	)and B(	63	);
	C	(	4051	)	<= A(	19	)and B(	63	);
	C	(	4052	)	<= A(	20	)and B(	63	);
	C	(	4053	)	<= A(	21	)and B(	63	);
	C	(	4054	)	<= A(	22	)and B(	63	);
	C	(	4055	)	<= A(	23	)and B(	63	);
	C	(	4056	)	<= A(	24	)and B(	63	);
	C	(	4057	)	<= A(	25	)and B(	63	);
	C	(	4058	)	<= A(	26	)and B(	63	);
	C	(	4059	)	<= A(	27	)and B(	63	);
	C	(	4060	)	<= A(	28	)and B(	63	);
	C	(	4061	)	<= A(	29	)and B(	63	);
	C	(	4062	)	<= A(	30	)and B(	63	);
	C	(	4063	)	<= A(	31	)and B(	63	);
	C	(	4064	)	<= A(	32	)and B(	63	);
	C	(	4065	)	<= A(	33	)and B(	63	);
	C	(	4066	)	<= A(	34	)and B(	63	);
	C	(	4067	)	<= A(	35	)and B(	63	);
	C	(	4068	)	<= A(	36	)and B(	63	);
	C	(	4069	)	<= A(	37	)and B(	63	);
	C	(	4070	)	<= A(	38	)and B(	63	);
	C	(	4071	)	<= A(	39	)and B(	63	);
	C	(	4072	)	<= A(	40	)and B(	63	);
	C	(	4073	)	<= A(	41	)and B(	63	);
	C	(	4074	)	<= A(	42	)and B(	63	);
	C	(	4075	)	<= A(	43	)and B(	63	);
	C	(	4076	)	<= A(	44	)and B(	63	);
	C	(	4077	)	<= A(	45	)and B(	63	);
	C	(	4078	)	<= A(	46	)and B(	63	);
	C	(	4079	)	<= A(	47	)and B(	63	);
	C	(	4080	)	<= A(	48	)and B(	63	);
	C	(	4081	)	<= A(	49	)and B(	63	);
	C	(	4082	)	<= A(	50	)and B(	63	);
	C	(	4083	)	<= A(	51	)and B(	63	);
	C	(	4084	)	<= A(	52	)and B(	63	);
	C	(	4085	)	<= A(	53	)and B(	63	);
	C	(	4086	)	<= A(	54	)and B(	63	);
	C	(	4087	)	<= A(	55	)and B(	63	);
	C	(	4088	)	<= A(	56	)and B(	63	);
	C	(	4089	)	<= A(	57	)and B(	63	);
	C	(	4090	)	<= A(	58	)and B(	63	);
	C	(	4091	)	<= A(	59	)and B(	63	);
	C	(	4092	)	<= A(	60	)and B(	63	);
	C	(	4093	)	<= A(	61	)and B(	63	);
	C	(	4094	)	<= A(	62	)and B(	63	);
	C	(	4095	)	<= A(	63	)and B(	63	);









--01-----------    
U0: Somador_Exato_1 PORT MAP(
   A => C(64),
   B => C(1),
   Cin => '0',
   Cout => Carry(0),
   S => R(1)
  );
 
U1: Somador_Exato_1 PORT MAP(
   A => C(65),
   B => C(2),
   Cin => Carry(0),
   Cout => Carry(1),
   S => E(0)
  );
 
U2: Somador_Exato_1 PORT MAP(
   A => C(66),
   B => C(3),
   Cin => Carry(1),
   Cout => Carry(2),
   S => E(1)
 );
 
U3: Somador_Exato_1 PORT MAP(
  A => C(67),
  B => C(4),
  Cin => Carry(2),
  Cout => Carry(3),
  S => E(2)
 );

 U4: Somador_Exato_1 PORT MAP(
  A => C(68),
  B => C(5),
  Cin => Carry(3),
  Cout => Carry(4),
  S => E(3)
 );
 
 U5: Somador_Exato_1 PORT MAP(
  A => C(69),
  B => C(6),
  Cin => Carry(4),
  Cout => Carry(5),
  S => E(4)
 ); 
 
 U6: Somador_Exato_1 PORT MAP(
  A => C(70),
  B => C(7),
  Cin => Carry(5),
  Cout => Carry(6),
  S => E(5)
 );  

 U7: Somador_Exato_1 PORT MAP(
  A => C(71),
  B => C(8),
  Cin => Carry(6),
  Cout => Carry(7),
  S => E(6)
 );  

 U8: Somador_Exato_1 PORT MAP(
  A => C(72),
  B => C(9),
  Cin => Carry(7),
  Cout => Carry(8),
  S => E(7)
 );  
 
 U9: Somador_Exato_1 PORT MAP(
  A => C(73),
  B => C(10),
  Cin => Carry(8),
  Cout => Carry(9),
  S => E(8)
 );  

 U10: Somador_Exato_1 PORT MAP(
  A => C(74),
  B => C(11),
  Cin => Carry(9),
  Cout => Carry(10),
  S => E(9)
 ); 
 
 U11: Somador_Exato_1 PORT MAP(
  A => C(75),
  B => C(12),
  Cin => Carry(10),
  Cout => Carry(11),
  S => E(10)
 ); 

 U12: Somador_Exato_1 PORT MAP(
  A => C(76),
  B => C(13),
  Cin => Carry(11),
  Cout => Carry(12),
  S => E(11)
 );

 U13: Somador_Exato_1 PORT MAP(
  A => C(77),
  B => C(14),
  Cin => Carry(12),
  Cout => Carry(13),
  S => E(12)
 ); 
 
 U14: Somador_Exato_1 PORT MAP(
  A => C(78),
  B => C(15),
  Cin => Carry(13),
  Cout => Carry(14),
  S => E(13)
 );
 
 U15: Somador_Exato_1 PORT MAP(
  A => C(79),
  B => C(16),
  Cin => Carry(14),
  Cout => Carry(15),
  S => E(14)
 );
 
 U16: Somador_Exato_1 PORT MAP(
  A => C(80),
  B => C(17),
  Cin => Carry(15),
  Cout => Carry(16),
  S => E(15)
 ); 
 
 U17: Somador_Exato_1 PORT MAP(
  A => C(81),
  B => C(18),
  Cin => Carry(16),
  Cout => Carry(17),
  S => E(16)
 );
 
 U18: Somador_Exato_1 PORT MAP(
  A => C(82),
  B => C(19),
  Cin => Carry(17),
  Cout => Carry(18),
  S => E(17)
 );
 
 U19: Somador_Exato_1 PORT MAP(
  A => C(83),
  B => C(20),
  Cin => Carry(18),
  Cout => Carry(19),
  S => E(18)
 ); 
 
 U20: Somador_Exato_1 PORT MAP(
  A => C(84),
  B => C(21),
  Cin => Carry(19),
  Cout => Carry(20),
  S => E(19)
 );

 U21: Somador_Exato_1 PORT MAP(
  A => C(85),
  B => C(22),
  Cin => Carry(20),
  Cout => Carry(21),
  S => E(20)
 ); 
 
 U22: Somador_Exato_1 PORT MAP(
  A => C(86),
  B => C(23),
  Cin => Carry(21),
  Cout => Carry(22),
  S => E(21)
 );
 
 U23: Somador_Exato_1 PORT MAP(
  A => C(87),
  B => C(24),
  Cin => Carry(22),
  Cout => Carry(23),
  S => E(22)
 );
 
 U24: Somador_Exato_1 PORT MAP(
  A => C(88),
  B => C(25),
  Cin => Carry(23),
  Cout => Carry(24),
  S => E(23)
 ); 
 
 U25: Somador_Exato_1 PORT MAP(
  A => C(89),
  B => C(26),
  Cin => Carry(24),
  Cout => Carry(25),
  S => E(24)
 );
 
 U26: Somador_Exato_1 PORT MAP(
  A => C(90),
  B => C(27),
  Cin => Carry(25),
  Cout => Carry(26),
  S => E(25)
 );
 
 U27: Somador_Exato_1 PORT MAP(
  A => C(91),
  B => C(28),
  Cin => Carry(26),
  Cout => Carry(27),
  S => E(26)
 ); 
 
 U28: Somador_Exato_1 PORT MAP(
  A => C(92),
  B => C(29),
  Cin => Carry(27),
  Cout => Carry(28),
  S => E(27)
 );

 U29: Somador_Exato_1 PORT MAP(
  A => C(93),
  B => C(30),
  Cin => Carry(28),
  Cout => Carry(29),
  S => E(28)
 ); 
 
 U30: Somador_Exato_1 PORT MAP(
  A => C(94),
  B => C(31),
  Cin => Carry(29),
  Cout => Carry(30),
  S => E(29)
 );
 
 U31: Somador_Exato_1 PORT MAP(
  A => C(95),
  B => C(32),
  Cin => Carry(30),
  Cout => Carry(31),
  S => E(30)
 );
 
 U32: Somador_Exato_1 PORT MAP(
  A => C(96),
  B => C(33),
  Cin => Carry(31),
  Cout => Carry(32),
  S => E(31)
 ); 
 
 U33: Somador_Exato_1 PORT MAP(
  A => C(97),
  B => C(34),
  Cin => Carry(32),
  Cout => Carry(33),
  S => E(32)
 );
 
 U34: Somador_Exato_1 PORT MAP(
  A => C(98),
  B => C(35),
  Cin => Carry(33),
  Cout => Carry(34),
  S => E(33)
 );
 
 U35: Somador_Exato_1 PORT MAP(
  A => C(99),
  B => C(36),
  Cin => Carry(34),
  Cout => Carry(35),
  S => E(34)
 ); 
 
 U36: Somador_Exato_1 PORT MAP(
  A => C(100),
  B => C(37),
  Cin => Carry(35),
  Cout => Carry(36),
  S => E(35)
 );

 U37: Somador_Exato_1 PORT MAP(
  A => C(101),
  B => C(38),
  Cin => Carry(36),
  Cout => Carry(37),
  S => E(36)
 ); 
 
 U38: Somador_Exato_1 PORT MAP(
  A => C(102),
  B => C(39),
  Cin => Carry(37),
  Cout => Carry(38),
  S => E(37)
 );
 
 U39: Somador_Exato_1 PORT MAP(
  A => C(103),
  B => C(40),
  Cin => Carry(38),
  Cout => Carry(39),
  S => E(38)
 );

 U40: Somador_Exato_1 PORT MAP(
  A => C(104),
  B => C(41),
  Cin => Carry(39),
  Cout => Carry(40),
  S => E(39)
 ); 
 
 U41: Somador_Exato_1 PORT MAP(
  A => C(105),
  B => C(42),
  Cin => Carry(40),
  Cout => Carry(41),
  S => E(40)
 );
 
 U42: Somador_Exato_1 PORT MAP(
  A => C(106),
  B => C(43),
  Cin => Carry(41),
  Cout => Carry(42),
  S => E(41)
 );
 
 U43: Somador_Exato_1 PORT MAP(
  A => C(107),
  B => C(44),
  Cin => Carry(42),
  Cout => Carry(43),
  S => E(42)
 ); 
 
 U44: Somador_Exato_1 PORT MAP(
  A => C(108),
  B => C(45),
  Cin => Carry(43),
  Cout => Carry(44),
  S => E(43)
 );

 U45: Somador_Exato_1 PORT MAP(
  A => C(109),
  B => C(46),
  Cin => Carry(44),
  Cout => Carry(45),
  S => E(44)
 ); 
 
 U46: Somador_Exato_1 PORT MAP(
  A => C(110),
  B => C(47),
  Cin => Carry(45),
  Cout => Carry(46),
  S => E(45)
 );
 
 U47: Somador_Exato_1 PORT MAP(
  A => C(111),
  B => C(48),
  Cin => Carry(46),
  Cout => Carry(47),
  S => E(46)
 );  
 
 U48: Somador_Exato_1 PORT MAP(
  A => C(112),
  B => C(49),
  Cin => Carry(47),
  Cout => Carry(48),
  S => E(47)
 ); 
 
 U49: Somador_Exato_1 PORT MAP(
  A => C(113),
  B => C(50),
  Cin => Carry(48),
  Cout => Carry(49),
  S => E(48)
 );
 
 U50: Somador_Exato_1 PORT MAP(
  A => C(114),
  B => C(51),
  Cin => Carry(49),
  Cout => Carry(50),
  S => E(49)
 );
 
 U51: Somador_Exato_1 PORT MAP(
  A => C(115),
  B => C(52),
  Cin => Carry(50),
  Cout => Carry(51),
  S => E(50)
 ); 
 
 U52: Somador_Exato_1 PORT MAP(
  A => C(116),
  B => C(53),
  Cin => Carry(51),
  Cout => Carry(52),
  S => E(51)
 );

 U53: Somador_Exato_1 PORT MAP(
  A => C(117),
  B => C(54),
  Cin => Carry(52),
  Cout => Carry(53),
  S => E(52)
 ); 
 
 U54: Somador_Exato_1 PORT MAP(
  A => C(118),
  B => C(55),
  Cin => Carry(53),
  Cout => Carry(54),
  S => E(53)
 );
 
 U55: Somador_Exato_1 PORT MAP(
  A => C(119),
  B => C(56),
  Cin => Carry(54),
  Cout => Carry(55),
  S => E(54)
 );

 U56: Somador_Exato_1 PORT MAP(
  A => C(120),
  B => E(57),
  Cin => Carry(55),
  Cout => Carry(56),
  S => E(55)
 ); 
 
 U57: Somador_Exato_1 PORT MAP(
  A => C(121),
  B => C(58),
  Cin => Carry(56),
  Cout => Carry(57),
  S => E(56)
 );
 
 U58: Somador_Exato_1 PORT MAP(
  A => C(122),
  B => C(59),
  Cin => Carry(57),
  Cout => Carry(58),
  S => E(57)
 );
 
 U59: Somador_Exato_1 PORT MAP(
  A => C(127),
  B => C(60),
  Cin => Carry(58),
  Cout => Carry(59),
  S => E(58)
 ); 
 
 U60: Somador_Exato_1 PORT MAP(
  A => C(124),
  B => C(61),
  Cin => Carry(59),
  Cout => Carry(60),
  S => E(59)
 );
 U61: Somador_Exato_1 PORT MAP(
  A => C(125),
  B => C(62),
  Cin => Carry(60),
  Cout => Carry(61),
  S => E(60)
 ); 
 
 U62: Somador_Exato_1 PORT MAP(
  A => C(126),
  B => C(63),
  Cin => Carry(61),
  Cout => Carry(62),
  S => E(61)
 );
 
 U63: Somador_Exato_1 PORT MAP(
  A => C(127),
  B => '0',
  Cin => Carry(62),
  Cout => Carry(63),
  S => E(62)
 );  

--2------
			
 U64	: Somador_Exato_1 PORT MAP(
	A=> C(	128	),
	B=>E(	0	),
	Cin=> '0'	,
	Cout=> Carry( 	64	),
	S=> R(	2	));
			
 U65	: Somador_Exato_1 PORT MAP(
	A=> C(	129	),
	B=>E(	1	),
	Cin=> Carry( 	64	),
	Cout=> Carry( 	65	),
	S=> E(	63	));
			
 U66	: Somador_Exato_1 PORT MAP(
	A=> C(	130	),
	B=>E(	2	),
	Cin=> Carry( 	65	),
	Cout=> Carry( 	66	),
	S=> E(	64	));
			
 U67	: Somador_Exato_1 PORT MAP(
	A=> C(	131	),
	B=>E(	3	),
	Cin=> Carry( 	66	),
	Cout=> Carry( 	67	),
	S=> E(	65	));
			
 U68	: Somador_Exato_1 PORT MAP(
	A=> C(	132	),
	B=>E(	4	),
	Cin=> Carry( 	67	),
	Cout=> Carry( 	68	),
	S=> E(	66	));
			
 U69	: Somador_Exato_1 PORT MAP(
	A=> C(	133	),
	B=>E(	5	),
	Cin=> Carry( 	68	),
	Cout=> Carry( 	69	),
	S=> E(	67	));
			
 U70	: Somador_Exato_1 PORT MAP(
	A=> C(	134	),
	B=>E(	6	),
	Cin=> Carry( 	69	),
	Cout=> Carry( 	70	),
	S=> E(	68	));
			
 U71	: Somador_Exato_1 PORT MAP(
	A=> C(	135	),
	B=>E(	7	),
	Cin=> Carry( 	70	),
	Cout=> Carry( 	71	),
	S=> E(	69	));
			
 U72	: Somador_Exato_1 PORT MAP(
	A=> C(	136	),
	B=>E(	8	),
	Cin=> Carry( 	71	),
	Cout=> Carry( 	72	),
	S=> E(	70	));
			
 U73	: Somador_Exato_1 PORT MAP(
	A=> C(	137	),
	B=>E(	9	),
	Cin=> Carry( 	72	),
	Cout=> Carry( 	73	),
	S=> E(	71	));
			
 U74	: Somador_Exato_1 PORT MAP(
	A=> C(	138	),
	B=>E(	10	),
	Cin=> Carry( 	73	),
	Cout=> Carry( 	74	),
	S=> E(	72	));
			
 U75	: Somador_Exato_1 PORT MAP(
	A=> C(	139	),
	B=>E(	11	),
	Cin=> Carry( 	74	),
	Cout=> Carry( 	75	),
	S=> E(	73	));
			
 U76	: Somador_Exato_1 PORT MAP(
	A=> C(	140	),
	B=>E(	12	),
	Cin=> Carry( 	75	),
	Cout=> Carry( 	76	),
	S=> E(	74	));
			
 U77	: Somador_Exato_1 PORT MAP(
	A=> C(	141	),
	B=>E(	13	),
	Cin=> Carry( 	76	),
	Cout=> Carry( 	77	),
	S=> E(	75	));
			
 U78	: Somador_Exato_1 PORT MAP(
	A=> C(	142	),
	B=>E(	14	),
	Cin=> Carry( 	77	),
	Cout=> Carry( 	78	),
	S=> E(	76	));
			
 U79	: Somador_Exato_1 PORT MAP(
	A=> C(	143	),
	B=>E(	15	),
	Cin=> Carry( 	78	),
	Cout=> Carry( 	79	),
	S=> E(	77	));
			
 U80	: Somador_Exato_1 PORT MAP(
	A=> C(	144	),
	B=>E(	16	),
	Cin=> Carry( 	79	),
	Cout=> Carry( 	80	),
	S=> E(	78	));
			
 U81	: Somador_Exato_1 PORT MAP(
	A=> C(	145	),
	B=>E(	17	),
	Cin=> Carry( 	80	),
	Cout=> Carry( 	81	),
	S=> E(	79	));
			
 U82	: Somador_Exato_1 PORT MAP(
	A=> C(	146	),
	B=>E(	18	),
	Cin=> Carry( 	81	),
	Cout=> Carry( 	82	),
	S=> E(	80	));
			
 U83	: Somador_Exato_1 PORT MAP(
	A=> C(	147	),
	B=>E(	19	),
	Cin=> Carry( 	82	),
	Cout=> Carry( 	83	),
	S=> E(	81	));
			
 U84	: Somador_Exato_1 PORT MAP(
	A=> C(	148	),
	B=>E(	20	),
	Cin=> Carry( 	83	),
	Cout=> Carry( 	84	),
	S=> E(	82	));
			
 U85	: Somador_Exato_1 PORT MAP(
	A=> C(	149	),
	B=>E(	21	),
	Cin=> Carry( 	84	),
	Cout=> Carry( 	85	),
	S=> E(	83	));
			
 U86	: Somador_Exato_1 PORT MAP(
	A=> C(	150	),
	B=>E(	22	),
	Cin=> Carry( 	85	),
	Cout=> Carry( 	86	),
	S=> E(	84	));
			
 U87	: Somador_Exato_1 PORT MAP(
	A=> C(	151	),
	B=>E(	23	),
	Cin=> Carry( 	86	),
	Cout=> Carry( 	87	),
	S=> E(	85	));
			
 U88	: Somador_Exato_1 PORT MAP(
	A=> C(	152	),
	B=>E(	24	),
	Cin=> Carry( 	87	),
	Cout=> Carry( 	88	),
	S=> E(	86	));
			
 U89	: Somador_Exato_1 PORT MAP(
	A=> C(	153	),
	B=>E(	25	),
	Cin=> Carry( 	88	),
	Cout=> Carry( 	89	),
	S=> E(	87	));
			
 U90	: Somador_Exato_1 PORT MAP(
	A=> C(	154	),
	B=>E(	26	),
	Cin=> Carry( 	89	),
	Cout=> Carry( 	90	),
	S=> E(	88	));
			
 U91	: Somador_Exato_1 PORT MAP(
	A=> C(	155	),
	B=>E(	27	),
	Cin=> Carry( 	90	),
	Cout=> Carry( 	91	),
	S=> E(	89	));
			
 U92	: Somador_Exato_1 PORT MAP(
	A=> C(	156	),
	B=>E(	28	),
	Cin=> Carry( 	91	),
	Cout=> Carry( 	92	),
	S=> E(	90	));
			
 U93	: Somador_Exato_1 PORT MAP(
	A=> C(	157	),
	B=>E(	29	),
	Cin=> Carry( 	92	),
	Cout=> Carry( 	93	),
	S=> E(	91	));
			
 U94	: Somador_Exato_1 PORT MAP(
	A=> C(	158	),
	B=>E(	30	),
	Cin=> Carry( 	93	),
	Cout=> Carry( 	94	),
	S=> E(	92	));
			
 U95	: Somador_Exato_1 PORT MAP(
	A=> C(	159	),
	B=>E(	31	),
	Cin=> Carry( 	94	),
	Cout=> Carry( 	95	),
	S=> E(	93	));
			
 U96	: Somador_Exato_1 PORT MAP(
	A=> C(	160	),
	B=>E(	32	),
	Cin=> Carry( 	95	),
	Cout=> Carry( 	96	),
	S=> E(	94	));
			
 U97	: Somador_Exato_1 PORT MAP(
	A=> C(	161	),
	B=>E(	33	),
	Cin=> Carry( 	96	),
	Cout=> Carry( 	97	),
	S=> E(	95	));
			
 U98	: Somador_Exato_1 PORT MAP(
	A=> C(	162	),
	B=>E(	34	),
	Cin=> Carry( 	97	),
	Cout=> Carry( 	98	),
	S=> E(	96	));
			
 U99	: Somador_Exato_1 PORT MAP(
	A=> C(	163	),
	B=>E(	35	),
	Cin=> Carry( 	98	),
	Cout=> Carry( 	99	),
	S=> E(	97	));
			
 U100	: Somador_Exato_1 PORT MAP(
	A=> C(	164	),
	B=>E(	36	),
	Cin=> Carry( 	99	),
	Cout=> Carry( 	100	),
	S=> E(	98	));
			
 U101	: Somador_Exato_1 PORT MAP(
	A=> C(	165	),
	B=>E(	37	),
	Cin=> Carry( 	100	),
	Cout=> Carry( 	101	),
	S=> E(	99	));
			
 U102	: Somador_Exato_1 PORT MAP(
	A=> C(	166	),
	B=>E(	38	),
	Cin=> Carry( 	101	),
	Cout=> Carry( 	102	),
	S=> E(	100	));
			
 U103	: Somador_Exato_1 PORT MAP(
	A=> C(	167	),
	B=>E(	39	),
	Cin=> Carry( 	102	),
	Cout=> Carry( 	103	),
	S=> E(	101	));
			
 U104	: Somador_Exato_1 PORT MAP(
	A=> C(	168	),
	B=>E(	40	),
	Cin=> Carry( 	103	),
	Cout=> Carry( 	104	),
	S=> E(	102	));
			
 U105	: Somador_Exato_1 PORT MAP(
	A=> C(	169	),
	B=>E(	41	),
	Cin=> Carry( 	104	),
	Cout=> Carry( 	105	),
	S=> E(	103	));
			
 U106	: Somador_Exato_1 PORT MAP(
	A=> C(	170	),
	B=>E(	42	),
	Cin=> Carry( 	105	),
	Cout=> Carry( 	106	),
	S=> E(	104	));
			
 U107	: Somador_Exato_1 PORT MAP(
	A=> C(	171	),
	B=>E(	43	),
	Cin=> Carry( 	106	),
	Cout=> Carry( 	107	),
	S=> E(	105	));
			
 U108	: Somador_Exato_1 PORT MAP(
	A=> C(	172	),
	B=> E(	44	),
	Cin=> Carry( 	107	),
	Cout=> Carry( 	108	),
	S=> E(	106	));
			
 U109	: Somador_Exato_1 PORT MAP(
	A=> C(	173	),
	B=> E(	45	),
	Cin=> Carry( 	108	),
	Cout=> Carry( 	109	),
	S=> E(	107	));
			
 U110	: Somador_Exato_1 PORT MAP(
	A=> C(	174	),
	B=> E(	46	),
	Cin=> Carry( 	109	),
	Cout=> Carry( 	110	),
	S=> E(	108	));
			
 U111	: Somador_Exato_1 PORT MAP(
	A=> C(	175	),
	B=> E(	47	),
	Cin=> Carry( 	110	),
	Cout=> Carry( 	111	),
	S=> E(	109	));
			
 U112	: Somador_Exato_1 PORT MAP(
	A=> C(	176	),
	B=> E(	48	),
	Cin=> Carry( 	111	),
	Cout=> Carry( 	112	),
	S=> E(	110	));
			
 U113	: Somador_Exato_1 PORT MAP(
	A=> C(	177	),
	B=> E(	49	),
	Cin=> Carry( 	112	),
	Cout=> Carry( 	113	),
	S=> E(	111	));
			
 U114	: Somador_Exato_1 PORT MAP(
	A=> C(	178	),
	B=> E(	50	),
	Cin=> Carry( 	113	),
	Cout=> Carry( 	114	),
	S=> E(	112	));
			
 U115	: Somador_Exato_1 PORT MAP(
	A=> C(	179	),
	B=> E(	51	),
	Cin=> Carry( 	114	),
	Cout=> Carry( 	115	),
	S=> E(	113	));
			
 U116	: Somador_Exato_1 PORT MAP(
	A=> C(	180	),
	B=> E(	52	),
	Cin=> Carry( 	115	),
	Cout=> Carry( 	116	),
	S=> E(	114	));
			
 U117	: Somador_Exato_1 PORT MAP(
	A=> C(	181	),
	B=> E(	53	),
	Cin=> Carry( 	116	),
	Cout=> Carry( 	117	),
	S=> E(	115	));
			
 U118	: Somador_Exato_1 PORT MAP(
	A=> C(	182	),
	B=>E(	54	),
	Cin=> Carry( 	117	),
	Cout=> Carry( 	118	),
	S=> E(	116	));
			
 U119	: Somador_Exato_1 PORT MAP(
	A=> C(	183	),
	B=> E(	55	),
	Cin=> Carry( 	118	),
	Cout=> Carry( 	119	),
	S=> E(	117	));
			
 U120	: Somador_Exato_1 PORT MAP(
	A=> C(	184	),
	B=> E(	56	),
	Cin=> Carry( 	119	),
	Cout=> Carry( 	120	),
	S=> E(	118	));
			
 U121	: Somador_Exato_1 PORT MAP(
	A=> C(	185	),
	B=> E(	57	),
	Cin=> Carry( 	120	),
	Cout=> Carry( 	121	),
	S=> E(	119	));
			
 U122	: Somador_Exato_1 PORT MAP(
	A=> C(	186	),
	B=> E(	58	),
	Cin=> Carry( 	121	),
	Cout=> Carry( 	122	),
	S=> E(	120	));
			
 U123	: Somador_Exato_1 PORT MAP(
	A=> C(	187	),
	B=> E(	59	),
	Cin=> Carry( 	122	),
	Cout=> Carry( 	123	),
	S=> E(	121	));
			
 U124	: Somador_Exato_1 PORT MAP(
	A=> C(	188	),
	B=> E(	60	),
	Cin=> Carry( 	123	),
	Cout=> Carry( 	124	),
	S=> E(	122	));
			
 U125	: Somador_Exato_1 PORT MAP(
	A=> C(	189	),
	B=> E(	61	),
	Cin=> Carry( 	124	),
	Cout=> Carry( 	125	),
	S=> E(	123	));
			
 U126	: Somador_Exato_1 PORT MAP(
	A=> C(	190	),
	B=> E(	62	),
	Cin=> Carry( 	125	),
	Cout=> Carry( 	126	),
	S=> E(	124	));
			
 U127	: Somador_Exato_1 PORT MAP(
	A => C(191),
	B => Carry(63),
	Cin => Carry(126),
	Cout => Carry(127),
	S=> E(	125	));
------3
			
 U128	: Somador_Exato_1 PORT MAP(
	A=> C(	192	),
	B=> E(	63	),
	Cin=> '0'	,
	Cout=> Carry( 	128	),
	S=> R(	3	));
			
 U129	: Somador_Exato_1 PORT MAP(
	A=> C(	193	),
	B=> E(	64	),
	Cin=> Carry( 	128	),
	Cout=> Carry( 	129	),
	S=> E(	126	));
			
 U130	: Somador_Exato_1 PORT MAP(
	A=> C(	194	),
	B=> E(	65	),
	Cin=> Carry( 	129	),
	Cout=> Carry( 	130	),
	S=> E(	127	));
			
 U131	: Somador_Exato_1 PORT MAP(
	A=> C(	195	),
	B=> E(	66	),
	Cin=> Carry( 	130	),
	Cout=> Carry( 	131	),
	S=> E(	128	));
			
 U132	: Somador_Exato_1 PORT MAP(
	A=> C(	196	),
	B=> E(	67	),
	Cin=> Carry( 	131	),
	Cout=> Carry( 	132	),
	S=> E(	129	));
			
 U133	: Somador_Exato_1 PORT MAP(
	A=> C(	197	),
	B=> E(	68	),
	Cin=> Carry( 	132	),
	Cout=> Carry( 	133	),
	S=> E(	130	));
			
 U134	: Somador_Exato_1 PORT MAP(
	A=> C(	198	),
	B=> E(	69	),
	Cin=> Carry( 	133	),
	Cout=> Carry( 	134	),
	S=> E(	131	));
			
 U135	: Somador_Exato_1 PORT MAP(
	A=> C(	199	),
	B=> E(	70	),
	Cin=> Carry( 	134	),
	Cout=> Carry( 	135	),
	S=> E(	132	));
			
 U136	: Somador_Exato_1 PORT MAP(
	A=> C(	200	),
	B=> E(	71	),
	Cin=> Carry( 	135	),
	Cout=> Carry( 	136	),
	S=> E(	133	));
			
 U137	: Somador_Exato_1 PORT MAP(
	A=> C(	201	),
	B=> E(	72	),
	Cin=> Carry( 	136	),
	Cout=> Carry( 	137	),
	S=> E(	134	));
			
 U138	: Somador_Exato_1 PORT MAP(
	A=> C(	202	),
	B=> E(	73	),
	Cin=> Carry( 	137	),
	Cout=> Carry( 	138	),
	S=> E(	135	));
			
 U139	: Somador_Exato_1 PORT MAP(
	A=> C(	203	),
	B=> E(	74	),
	Cin=> Carry( 	138	),
	Cout=> Carry( 	139	),
	S=> E(	136	));
			
 U140	: Somador_Exato_1 PORT MAP(
	A=> C(	204	),
	B=> E(	75	),
	Cin=> Carry( 	139	),
	Cout=> Carry( 	140	),
	S=> E(	137	));
			
 U141	: Somador_Exato_1 PORT MAP(
	A=> C(	205	),
	B=> E(	76	),
	Cin=> Carry( 	140	),
	Cout=> Carry( 	141	),
	S=> E(	138	));
			
 U142	: Somador_Exato_1 PORT MAP(
	A=> C(	206	),
	B=> E(	77	),
	Cin=> Carry( 	141	),
	Cout=> Carry( 	142	),
	S=> E(	139	));
			
 U143	: Somador_Exato_1 PORT MAP(
	A=> C(	207	),
	B=> E(	78	),
	Cin=> Carry( 	142	),
	Cout=> Carry( 	143	),
	S=> E(	140	));
			
 U144	: Somador_Exato_1 PORT MAP(
	A=> C(	208	),
	B=> E(	79	),
	Cin=> Carry( 	143	),
	Cout=> Carry( 	144	),
	S=> E(	141	));
			
 U145	: Somador_Exato_1 PORT MAP(
	A=> C(	209	),
	B=> E(	80	),
	Cin=> Carry( 	144	),
	Cout=> Carry( 	145	),
	S=> E(	142	));
			
 U146	: Somador_Exato_1 PORT MAP(
	A=> C(	210	),
	B=> E(	81	),
	Cin=> Carry( 	145	),
	Cout=> Carry( 	146	),
	S=> E(	143	));
			
 U147	: Somador_Exato_1 PORT MAP(
	A=> C(	211	),
	B=> E(	82	),
	Cin=> Carry( 	146	),
	Cout=> Carry( 	147	),
	S=> E(	144	));
			
 U148	: Somador_Exato_1 PORT MAP(
	A=> C(	212	),
	B=> E(	83	),
	Cin=> Carry( 	147	),
	Cout=> Carry( 	148	),
	S=> E(	145	));
			
 U149	: Somador_Exato_1 PORT MAP(
	A=> C(	213	),
	B=> E(	84	),
	Cin=> Carry( 	148	),
	Cout=> Carry( 	149	),
	S=> E(	146	));
			
 U150	: Somador_Exato_1 PORT MAP(
	A=> C(	214	),
	B=> E(	85	),
	Cin=> Carry( 	149	),
	Cout=> Carry( 	150	),
	S=> E(	147	));
			
 U151	: Somador_Exato_1 PORT MAP(
	A=> C(	215	),
	B=> E(	86	),
	Cin=> Carry( 	150	),
	Cout=> Carry( 	151	),
	S=> E(	148	));
			
 U152	: Somador_Exato_1 PORT MAP(
	A=> C(	216	),
	B=> E(	87	),
	Cin=> Carry( 	151	),
	Cout=> Carry( 	152	),
	S=> E(	149	));
			
 U153	: Somador_Exato_1 PORT MAP(
	A=> C(	217	),
	B=> E(	88	),
	Cin=> Carry( 	152	),
	Cout=> Carry( 	153	),
	S=> E(	150	));
			
 U154	: Somador_Exato_1 PORT MAP(
	A=> C(	218	),
	B=> E(	89	),
	Cin=> Carry( 	153	),
	Cout=> Carry( 	154	),
	S=> E(	151	));
			
 U155	: Somador_Exato_1 PORT MAP(
	A=> C(	219	),
	B=> E(	90	),
	Cin=> Carry( 	154	),
	Cout=> Carry( 	155	),
	S=> E(	152	));
			
 U156	: Somador_Exato_1 PORT MAP(
	A=> C(	220	),
	B=> E(	91	),
	Cin=> Carry( 	155	),
	Cout=> Carry( 	156	),
	S=> E(	153	));
			
 U157	: Somador_Exato_1 PORT MAP(
	A=> C(	221	),
	B=> E(	92	),
	Cin=> Carry( 	156	),
	Cout=> Carry( 	157	),
	S=> E(	154	));
			
 U158	: Somador_Exato_1 PORT MAP(
	A=> C(	222	),
	B=> E(	93	),
	Cin=> Carry( 	157	),
	Cout=> Carry( 	158	),
	S=> E(	155	));
			
 U159	: Somador_Exato_1 PORT MAP(
	A=> C(	223	),
	B=> E(	94	),
	Cin=> Carry( 	158	),
	Cout=> Carry( 	159	),
	S=> E(	156	));
			
 U160	: Somador_Exato_1 PORT MAP(
	A=> C(	224	),
	B=> E(	95	),
	Cin=> Carry( 	159	),
	Cout=> Carry( 	160	),
	S=> E(	157	));
			
 U161	: Somador_Exato_1 PORT MAP(
	A=> C(	225	),
	B=> E(	96	),
	Cin=> Carry( 	160	),
	Cout=> Carry( 	161	),
	S=> E(	158	));
			
 U162	: Somador_Exato_1 PORT MAP(
	A=> C(	226	),
	B=> E(	97	),
	Cin=> Carry( 	161	),
	Cout=> Carry( 	162	),
	S=> E(	159	));
			
 U163	: Somador_Exato_1 PORT MAP(
	A=> C(	227	),
	B=> E(	98	),
	Cin=> Carry( 	162	),
	Cout=> Carry( 	163	),
	S=> E(	160	));
			
 U164	: Somador_Exato_1 PORT MAP(
	A=> C(	228	),
	B=> E(	99	),
	Cin=> Carry( 	163	),
	Cout=> Carry( 	164	),
	S=> E(	161	));
			
 U165	: Somador_Exato_1 PORT MAP(
	A=> C(	229	),
	B=> E(	100	),
	Cin=> Carry( 	164	),
	Cout=> Carry( 	165	),
	S=> E(	162	));
			
 U166	: Somador_Exato_1 PORT MAP(
	A=> C(	230	),
	B=> E(	101	),
	Cin=> Carry( 	165	),
	Cout=> Carry( 	166	),
	S=> E(	163	));
			
 U167	: Somador_Exato_1 PORT MAP(
	A=> C(	231	),
	B=> E(	102	),
	Cin=> Carry( 	166	),
	Cout=> Carry( 	167	),
	S=> E(	164	));
			
 U168	: Somador_Exato_1 PORT MAP(
	A=> C(	232	),
	B=> E(	103	),
	Cin=> Carry( 	167	),
	Cout=> Carry( 	168	),
	S=> E(	165	));
			
 U169	: Somador_Exato_1 PORT MAP(
	A=> C(	233	),
	B=> E(	104	),
	Cin=> Carry( 	168	),
	Cout=> Carry( 	169	),
	S=> E(	166	));
			
 U170	: Somador_Exato_1 PORT MAP(
	A=> C(	234	),
	B=> E(	105	),
	Cin=> Carry( 	169	),
	Cout=> Carry( 	170	),
	S=> E(	167	));
			
 U171	: Somador_Exato_1 PORT MAP(
	A=> C(	235	),
	B=> E(	106	),
	Cin=> Carry( 	170	),
	Cout=> Carry( 	171	),
	S=> E(	168	));
			
 U172	: Somador_Exato_1 PORT MAP(
	A=> C(	236	),
	B=> E(	107	),
	Cin=> Carry( 	171	),
	Cout=> Carry( 	172	),
	S=> E(	169	));
			
 U173	: Somador_Exato_1 PORT MAP(
	A=> C(	237	),
	B=> E(	108	),
	Cin=> Carry( 	172	),
	Cout=> Carry( 	173	),
	S=> E(	170	));
			
 U174	: Somador_Exato_1 PORT MAP(
	A=> C(	238	),
	B=> E(	109	),
	Cin=> Carry( 	173	),
	Cout=> Carry( 	174	),
	S=> E(	171	));
			
 U175	: Somador_Exato_1 PORT MAP(
	A=> C(	239	),
	B=> E(	110	),
	Cin=> Carry( 	174	),
	Cout=> Carry( 	175	),
	S=> E(	172	));
			
 U176	: Somador_Exato_1 PORT MAP(
	A=> C(	240	),
	B=> E(	111	),
	Cin=> Carry( 	175	),
	Cout=> Carry( 	176	),
	S=> E(	173	));
			
 U177	: Somador_Exato_1 PORT MAP(
	A=> C(	241	),
	B=> E(	112	),
	Cin=> Carry( 	176	),
	Cout=> Carry( 	177	),
	S=> E(	174	));
			
 U178	: Somador_Exato_1 PORT MAP(
	A=> C(	242	),
	B=> E(	113	),
	Cin=> Carry( 	177	),
	Cout=> Carry( 	178	),
	S=> E(	175	));
			
 U179	: Somador_Exato_1 PORT MAP(
	A=> C(	243	),
	B=> E(	114	),
	Cin=> Carry( 	178	),
	Cout=> Carry( 	179	),
	S=> E(	176	));
			
 U180	: Somador_Exato_1 PORT MAP(
	A=> C(	244	),
	B=> E(	115	),
	Cin=> Carry( 	179	),
	Cout=> Carry( 	180	),
	S=> E(	177	));
			
 U181	: Somador_Exato_1 PORT MAP(
	A=> C(	245	),
	B=> E(	116	),
	Cin=> Carry( 	180	),
	Cout=> Carry( 	181	),
	S=> E(	178	));
			
 U182	: Somador_Exato_1 PORT MAP(
	A=> C(	246	),
	B=> E(	117	),
	Cin=> Carry( 	181	),
	Cout=> Carry( 	182	),
	S=> E(	179	));
			
 U183	: Somador_Exato_1 PORT MAP(
	A=> C(	247	),
	B=> E(	118	),
	Cin=> Carry( 	182	),
	Cout=> Carry( 	183	),
	S=> E(	180	));
			
 U184	: Somador_Exato_1 PORT MAP(
	A=> C(	248	),
	B=> E(	119	),
	Cin=> Carry( 	183	),
	Cout=> Carry( 	184	),
	S=> E(	181	));
			
 U185	: Somador_Exato_1 PORT MAP(
	A=> C(	249	),
	B=> E(	120	),
	Cin=> Carry( 	184	),
	Cout=> Carry( 	185	),
	S=> E(	182	));
			
 U186	: Somador_Exato_1 PORT MAP(
	A=> C(	250	),
	B=> E(	121	),
	Cin=> Carry( 	185	),
	Cout=> Carry( 	186	),
	S=> E(	183	));
			
 U187	: Somador_Exato_1 PORT MAP(
	A=> C(	251	),
	B=> E(	122	),
	Cin=> Carry( 	186	),
	Cout=> Carry( 	187	),
	S=> E(	184	));
			
 U188	: Somador_Exato_1 PORT MAP(
	A=> C(	252	),
	B=> E(	123	),
	Cin=> Carry( 	187	),
	Cout=> Carry( 	188	),
	S=> E(	185	));
			
 U189	: Somador_Exato_1 PORT MAP(
	A=> C(	253	),
	B=> E(	124	),
	Cin=> Carry( 	188	),
	Cout=> Carry( 	189	),
	S=> E(	186	));
			
 U190	: Somador_Exato_1 PORT MAP(
	A=> C(	254	),
	B=> E(	125	),
	Cin=> Carry( 	189	),
	Cout=> Carry( 	190	),
	S=> E(	187	));
			
 U191	: Somador_Exato_1 PORT MAP(
	A => C(255),
	B => Carry(127),
	Cin => Carry(190),
	Cout => Carry(191),
	S => E(188));
---4
				
 U192	: Somador_Exato_1 PORT MAP(	
	A=> C(	256	),	
	B=> E(	126	),	
	Cin=> '0'	,	
	Cout=> Carry( 	192	),	
	S=> R(	4	));	
				
 U193	: Somador_Exato_1 PORT MAP(	
	A=> C(	257	),	
	B=> E(	127	),	
	Cin=> Carry( 	192	),	
	Cout=> Carry( 	193	),	
	S=> E(	189	));	
				
 U194	: Somador_Exato_1 PORT MAP(	
	A=> C(	258	),	
	B=> E(	128	),	
	Cin=> Carry( 	193	),	
	Cout=> Carry( 	194	),	
	S=> E(	190	));	
				
 U195	: Somador_Exato_1 PORT MAP(	
	A=> C(	259	),	
	B=> E(	129	),	
	Cin=> Carry( 	194	),	
	Cout=> Carry( 	195	),	
	S=> E(	191	));	
				
 U196	: Somador_Exato_1 PORT MAP(	
	A=> C(	260	),	
	B=> E(	130	),	
	Cin=> Carry( 	195	),	
	Cout=> Carry( 	196	),	
	S=> E(	192	));	
				
 U197	: Somador_Exato_1 PORT MAP(	
	A=> C(	261	),	
	B=> E(	131	),	
	Cin=> Carry( 	196	),	
	Cout=> Carry( 	197	),	
	S=> E(	193	));	
				
 U198	: Somador_Exato_1 PORT MAP(	
	A=> C(	262	),	
	B=> E(	132	),	
	Cin=> Carry( 	197	),	
	Cout=> Carry( 	198	),	
	S=> E(	194	));	
				
 U199	: Somador_Exato_1 PORT MAP(	
	A=> C(	263	),	
	B=> E(	133	),	
	Cin=> Carry( 	198	),	
	Cout=> Carry( 	199	),	
	S=> E(	195	));	
				
 U200	: Somador_Exato_1 PORT MAP(	
	A=> C(	264	),	
	B=> E(	134	),	
	Cin=> Carry( 	199	),	
	Cout=> Carry( 	200	),	
	S=> E(	196	));	
				
 U201	: Somador_Exato_1 PORT MAP(	
	A=> C(	265	),	
	B=> E(	135	),	
	Cin=> Carry( 	200	),	
	Cout=> Carry( 	201	),	
	S=> E(	197	));	
				
 U202	: Somador_Exato_1 PORT MAP(	
	A=> C(	266	),	
	B=> E(	136	),	
	Cin=> Carry( 	201	),	
	Cout=> Carry( 	202	),	
	S=> E(	198	));	
				
 U203	: Somador_Exato_1 PORT MAP(	
	A=> C(	267	),	
	B=> E(	137	),	
	Cin=> Carry( 	202	),	
	Cout=> Carry( 	203	),	
	S=> E(	199	));	
				
 U204	: Somador_Exato_1 PORT MAP(	
	A=> C(	268	),	
	B=> E(	138	),	
	Cin=> Carry( 	203	),	
	Cout=> Carry( 	204	),	
	S=> E(	200	));	
				
 U205	: Somador_Exato_1 PORT MAP(	
	A=> C(	269	),	
	B=> E(	139	),	
	Cin=> Carry( 	204	),	
	Cout=> Carry( 	205	),	
	S=> E(	201	));	
				
 U206	: Somador_Exato_1 PORT MAP(	
	A=> C(	270	),	
	B=> E(	140	),	
	Cin=> Carry( 	205	),	
	Cout=> Carry( 	206	),	
	S=> E(	202	));	
				
 U207	: Somador_Exato_1 PORT MAP(	
	A=> C(	271	),	
	B=> E(	141	),	
	Cin=> Carry( 	206	),	
	Cout=> Carry( 	207	),	
	S=> E(	203	));	
				
 U208	: Somador_Exato_1 PORT MAP(	
	A=> C(	272	),	
	B=> E(	142	),	
	Cin=> Carry( 	207	),	
	Cout=> Carry( 	208	),	
	S=> E(	204	));	
				
 U209	: Somador_Exato_1 PORT MAP(	
	A=> C(	273	),	
	B=> E(	143	),	
	Cin=> Carry( 	208	),	
	Cout=> Carry( 	209	),	
	S=> E(	205	));	
				
 U210	: Somador_Exato_1 PORT MAP(	
	A=> C(	274	),	
	B=> E(	144	),	
	Cin=> Carry( 	209	),	
	Cout=> Carry( 	210	),	
	S=> E(	206	));	
				
 U211	: Somador_Exato_1 PORT MAP(	
	A=> C(	275	),	
	B=> E(	145	),	
	Cin=> Carry( 	210	),	
	Cout=> Carry( 	211	),	
	S=> E(	207	));	
				
 U212	: Somador_Exato_1 PORT MAP(	
	A=> C(	276	),	
	B=> E(	146	),	
	Cin=> Carry( 	211	),	
	Cout=> Carry( 	212	),	
	S=> E(	208	));	
				
 U213	: Somador_Exato_1 PORT MAP(	
	A=> C(	277	),	
	B=> E(	147	),	
	Cin=> Carry( 	212	),	
	Cout=> Carry( 	213	),	
	S=> E(	209	));	
				
 U214	: Somador_Exato_1 PORT MAP(	
	A=> C(	278	),	
	B=> E(	148	),	
	Cin=> Carry( 	213	),	
	Cout=> Carry( 	214	),	
	S=> E(	210	));	
				
 U215	: Somador_Exato_1 PORT MAP(	
	A=> C(	279	),	
	B=> E(	149	),	
	Cin=> Carry( 	214	),	
	Cout=> Carry( 	215	),	
	S=> E(	211	));	
				
 U216	: Somador_Exato_1 PORT MAP(	
	A=> C(	280	),	
	B=> E(	150	),	
	Cin=> Carry( 	215	),	
	Cout=> Carry( 	216	),	
	S=> E(	212	));	
				
 U217	: Somador_Exato_1 PORT MAP(	
	A=> C(	281	),	
	B=> E(	151	),	
	Cin=> Carry( 	216	),	
	Cout=> Carry( 	217	),	
	S=> E(	213	));	
				
 U218	: Somador_Exato_1 PORT MAP(	
	A=> C(	282	),	
	B=> E(	152	),	
	Cin=> Carry( 	217	),	
	Cout=> Carry( 	218	),	
	S=> E(	214	));	
				
 U219	: Somador_Exato_1 PORT MAP(	
	A=> C(	283	),	
	B=> E(	153	),	
	Cin=> Carry( 	218	),	
	Cout=> Carry( 	219	),	
	S=> E(	215	));	
				
 U220	: Somador_Exato_1 PORT MAP(	
	A=> C(	284	),	
	B=> E(	154	),	
	Cin=> Carry( 	219	),	
	Cout=> Carry( 	220	),	
	S=> E(	216	));	
				
 U221	: Somador_Exato_1 PORT MAP(	
	A=> C(	285	),	
	B=> E(	155	),	
	Cin=> Carry( 	220	),	
	Cout=> Carry( 	221	),	
	S=> E(	217	));	
				
 U222	: Somador_Exato_1 PORT MAP(	
	A=> C(	286	),	
	B=> E(	156	),	
	Cin=> Carry( 	221	),	
	Cout=> Carry( 	222	),	
	S=> E(	218	));	
				
 U223	: Somador_Exato_1 PORT MAP(	
	A=> C(	287	),	
	B=> E(	157	),	
	Cin=> Carry( 	222	),	
	Cout=> Carry( 	223	),	
	S=> E(	219	));	
				
 U224	: Somador_Exato_1 PORT MAP(	
	A=> C(	288	),	
	B=> E(	158	),	
	Cin=> Carry( 	223	),	
	Cout=> Carry( 	224	),	
	S=> E(	220	));	
				
 U225	: Somador_Exato_1 PORT MAP(	
	A=> C(	289	),	
	B=> E(	159	),	
	Cin=> Carry( 	224	),	
	Cout=> Carry( 	225	),	
	S=> E(	221	));	
				
 U226	: Somador_Exato_1 PORT MAP(	
	A=> C(	290	),	
	B=> E(	160	),	
	Cin=> Carry( 	225	),	
	Cout=> Carry( 	226	),	
	S=> E(	222	));	
				
 U227	: Somador_Exato_1 PORT MAP(	
	A=> C(	291	),	
	B=> E(	161	),	
	Cin=> Carry( 	226	),	
	Cout=> Carry( 	227	),	
	S=> E(	223	));	
				
 U228	: Somador_Exato_1 PORT MAP(	
	A=> C(	292	),	
	B=> E(	162	),	
	Cin=> Carry( 	227	),	
	Cout=> Carry( 	228	),	
	S=> E(	224	));	
				
 U229	: Somador_Exato_1 PORT MAP(	
	A=> C(	293	),	
	B=> E(	163	),	
	Cin=> Carry( 	228	),	
	Cout=> Carry( 	229	),	
	S=> E(	225	));	
				
 U230	: Somador_Exato_1 PORT MAP(	
	A=> C(	294	),	
	B=> E(	164	),	
	Cin=> Carry( 	229	),	
	Cout=> Carry( 	230	),	
	S=> E(	226	));	
				
 U231	: Somador_Exato_1 PORT MAP(	
	A=> C(	295	),	
	B=> E(	165	),	
	Cin=> Carry( 	230	),	
	Cout=> Carry( 	231	),	
	S=> E(	227	));	
				
 U232	: Somador_Exato_1 PORT MAP(	
	A=> C(	296	),	
	B=> E(	166	),	
	Cin=> Carry( 	231	),	
	Cout=> Carry( 	232	),	
	S=> E(	228	));	
				
 U233	: Somador_Exato_1 PORT MAP(	
	A=> C(	297	),	
	B=> E(	167	),	
	Cin=> Carry( 	232	),	
	Cout=> Carry( 	233	),	
	S=> E(	229	));	
				
 U234	: Somador_Exato_1 PORT MAP(	
	A=> C(	298	),	
	B=> E(	168	),	
	Cin=> Carry( 	233	),	
	Cout=> Carry( 	234	),	
	S=> E(	230	));	
				
 U235	: Somador_Exato_1 PORT MAP(	
	A=> C(	299	),	
	B=> E(	169	),	
	Cin=> Carry( 	234	),	
	Cout=> Carry( 	235	),	
	S=> E(	231	));	
				
 U236	: Somador_Exato_1 PORT MAP(	
	A=> C(	300	),	
	B=> E(	170	),	
	Cin=> Carry( 	235	),	
	Cout=> Carry( 	236	),	
	S=> E(	232	));	
				
 U237	: Somador_Exato_1 PORT MAP(	
	A=> C(	301	),	
	B=> E(	171	),	
	Cin=> Carry( 	236	),	
	Cout=> Carry( 	237	),	
	S=> E(	233	));	
				
 U238	: Somador_Exato_1 PORT MAP(	
	A=> C(	302	),	
	B=> E(	172	),	
	Cin=> Carry( 	237	),	
	Cout=> Carry( 	238	),	
	S=> E(	234	));	
				
 U239	: Somador_Exato_1 PORT MAP(	
	A=> C(	303	),	
	B=> E(	173	),	
	Cin=> Carry( 	238	),	
	Cout=> Carry( 	239	),	
	S=> E(	235	));	
				
 U240	: Somador_Exato_1 PORT MAP(	
	A=> C(	304	),	
	B=> E(	174	),	
	Cin=> Carry( 	239	),	
	Cout=> Carry( 	240	),	
	S=> E(	236	));	
				
 U241	: Somador_Exato_1 PORT MAP(	
	A=> C(	305	),	
	B=> E(	175	),	
	Cin=> Carry( 	240	),	
	Cout=> Carry( 	241	),	
	S=> E(	237	));	
				
 U242	: Somador_Exato_1 PORT MAP(	
	A=> C(	306	),	
	B=> E(	176	),	
	Cin=> Carry( 	241	),	
	Cout=> Carry( 	242	),	
	S=> E(	238	));	
				
 U243	: Somador_Exato_1 PORT MAP(	
	A=> C(	307	),	
	B=> E(	177	),	
	Cin=> Carry( 	242	),	
	Cout=> Carry( 	243	),	
	S=> E(	239	));	
				
 U244	: Somador_Exato_1 PORT MAP(	
	A=> C(	308	),	
	B=> E(	178	),	
	Cin=> Carry( 	243	),	
	Cout=> Carry( 	244	),	
	S=> E(	240	));	
				
 U245	: Somador_Exato_1 PORT MAP(	
	A=> C(	309	),	
	B=> E(	179	),	
	Cin=> Carry( 	244	),	
	Cout=> Carry( 	245	),	
	S=> E(	241	));	
				
 U246	: Somador_Exato_1 PORT MAP(	
	A=> C(	310	),	
	B=> E(	180	),	
	Cin=> Carry( 	245	),	
	Cout=> Carry( 	246	),	
	S=> E(	242	));	
				
 U247	: Somador_Exato_1 PORT MAP(	
	A=> C(	311	),	
	B=> E(	181	),	
	Cin=> Carry( 	246	),	
	Cout=> Carry( 	247	),	
	S=> E(	243	));	
				
 U248	: Somador_Exato_1 PORT MAP(	
	A=> C(	312	),	
	B=> E(	182	),	
	Cin=> Carry( 	247	),	
	Cout=> Carry( 	248	),	
	S=> E(	244	));	
				
 U249	: Somador_Exato_1 PORT MAP(	
	A=> C(	313	),	
	B=> E(	183	),	
	Cin=> Carry( 	248	),	
	Cout=> Carry( 	249	),	
	S=> E(	245	));	
				
 U250	: Somador_Exato_1 PORT MAP(	
	A=> C(	314	),	
	B=> E(	184	),	
	Cin=> Carry( 	249	),	
	Cout=> Carry( 	250	),	
	S=> E(	246	));	
				
 U251	: Somador_Exato_1 PORT MAP(	
	A=> C(	315	),	
	B=> E(	185	),	
	Cin=> Carry( 	250	),	
	Cout=> Carry( 	251	),	
	S=> E(	247	));	
				
 U252	: Somador_Exato_1 PORT MAP(	
	A=> C(	316	),	
	B=> E(	186	),	
	Cin=> Carry( 	251	),	
	Cout=> Carry( 	252	),	
	S=> E(	248	));	
				
 U253	: Somador_Exato_1 PORT MAP(	
	A=> C(	317	),	
	B=> E(	187	),	
	Cin=> Carry( 	252	),	
	Cout=> Carry( 	253	),	
	S=> E(	249	));	
				
 U254	: Somador_Exato_1 PORT MAP(	
	A=> C(	318	),	
	B=> E(	188	),	
	Cin=> Carry( 	253	),	
	Cout=> Carry( 	254	),	
	S=> E(	250	));	
				
 U255	: Somador_Exato_1 PORT MAP(	
	A => C(319),	
	B => Carry(191),	
	Cin => Carry(254),	
	Cout => Carry(255),	
	S => E(	251	));	
---5
			
 U256	: Somador_Exato_1 PORT MAP(
	A=> C(	320	),
	B=> E(	189	),
	Cin=> '0'	,
	Cout=> Carry( 	256	),
	S=> R(	5	));
			
 U257	: Somador_Exato_1 PORT MAP(
	A=> C(	321	),
	B=> E(	190	),
	Cin=> Carry( 	256	),
	Cout=> Carry( 	257	),
	S=> E(	252	));
			
 U258	: Somador_Exato_1 PORT MAP(
	A=> C(	322	),
	B=> E(	191	),
	Cin=> Carry( 	257	),
	Cout=> Carry( 	258	),
	S=> E(	253	));
			
 U259	: Somador_Exato_1 PORT MAP(
	A=> C(	323	),
	B=> E(	192	),
	Cin=> Carry( 	258	),
	Cout=> Carry( 	259	),
	S=> E(	254	));
			
 U260	: Somador_Exato_1 PORT MAP(
	A=> C(	324	),
	B=> E(	193	),
	Cin=> Carry( 	259	),
	Cout=> Carry( 	260	),
	S=> E(	255	));
			
 U261	: Somador_Exato_1 PORT MAP(
	A=> C(	325	),
	B=> E(	194	),
	Cin=> Carry( 	260	),
	Cout=> Carry( 	261	),
	S=> E(	256	));
			
 U262	: Somador_Exato_1 PORT MAP(
	A=> C(	326	),
	B=> E(	195	),
	Cin=> Carry( 	261	),
	Cout=> Carry( 	262	),
	S=> E(	257	));
			
 U263	: Somador_Exato_1 PORT MAP(
	A=> C(	327	),
	B=> E(	196	),
	Cin=> Carry( 	262	),
	Cout=> Carry( 	263	),
	S=> E(	258	));
			
 U264	: Somador_Exato_1 PORT MAP(
	A=> C(	328	),
	B=> E(	197	),
	Cin=> Carry( 	263	),
	Cout=> Carry( 	264	),
	S=> E(	259	));
			
 U265	: Somador_Exato_1 PORT MAP(
	A=> C(	329	),
	B=> E(	198	),
	Cin=> Carry( 	264	),
	Cout=> Carry( 	265	),
	S=> E(	260	));
			
 U266	: Somador_Exato_1 PORT MAP(
	A=> C(	330	),
	B=> E(	199	),
	Cin=> Carry( 	265	),
	Cout=> Carry( 	266	),
	S=> E(	261	));
			
 U267	: Somador_Exato_1 PORT MAP(
	A=> C(	331	),
	B=> E(	200	),
	Cin=> Carry( 	266	),
	Cout=> Carry( 	267	),
	S=> E(	262	));
			
 U268	: Somador_Exato_1 PORT MAP(
	A=> C(	332	),
	B=> E(	201	),
	Cin=> Carry( 	267	),
	Cout=> Carry( 	268	),
	S=> E(	263	));
			
 U269	: Somador_Exato_1 PORT MAP(
	A=> C(	333	),
	B=> E(	202	),
	Cin=> Carry( 	268	),
	Cout=> Carry( 	269	),
	S=> E(	264	));
			
 U270	: Somador_Exato_1 PORT MAP(
	A=> C(	334	),
	B=> E(	203	),
	Cin=> Carry( 	269	),
	Cout=> Carry( 	270	),
	S=> E(	265	));
			
 U271	: Somador_Exato_1 PORT MAP(
	A=> C(	335	),
	B=> E(	204	),
	Cin=> Carry( 	270	),
	Cout=> Carry( 	271	),
	S=> E(	266	));
			
 U272	: Somador_Exato_1 PORT MAP(
	A=> C(	336	),
	B=> E(	205	),
	Cin=> Carry( 	271	),
	Cout=> Carry( 	272	),
	S=> E(	267	));
			
 U273	: Somador_Exato_1 PORT MAP(
	A=> C(	337	),
	B=> E(	206	),
	Cin=> Carry( 	272	),
	Cout=> Carry( 	273	),
	S=> E(	268	));
			
 U274	: Somador_Exato_1 PORT MAP(
	A=> C(	338	),
	B=> E(	207	),
	Cin=> Carry( 	273	),
	Cout=> Carry( 	274	),
	S=> E(	269	));
			
 U275	: Somador_Exato_1 PORT MAP(
	A=> C(	339	),
	B=> E(	208	),
	Cin=> Carry( 	274	),
	Cout=> Carry( 	275	),
	S=> E(	270	));
			
 U276	: Somador_Exato_1 PORT MAP(
	A=> C(	340	),
	B=> E(	209	),
	Cin=> Carry( 	275	),
	Cout=> Carry( 	276	),
	S=> E(	271	));
			
 U277	: Somador_Exato_1 PORT MAP(
	A=> C(	341	),
	B=> E(	210	),
	Cin=> Carry( 	276	),
	Cout=> Carry( 	277	),
	S=> E(	272	));
			
 U278	: Somador_Exato_1 PORT MAP(
	A=> C(	342	),
	B=> E(	211	),
	Cin=> Carry( 	277	),
	Cout=> Carry( 	278	),
	S=> E(	273	));
			
 U279	: Somador_Exato_1 PORT MAP(
	A=> C(	343	),
	B=> E(	212	),
	Cin=> Carry( 	278	),
	Cout=> Carry( 	279	),
	S=> E(	274	));
			
 U280	: Somador_Exato_1 PORT MAP(
	A=> C(	344	),
	B=> E(	213	),
	Cin=> Carry( 	279	),
	Cout=> Carry( 	280	),
	S=> E(	275	));
			
 U281	: Somador_Exato_1 PORT MAP(
	A=> C(	345	),
	B=> E(	214	),
	Cin=> Carry( 	280	),
	Cout=> Carry( 	281	),
	S=> E(	276	));
			
 U282	: Somador_Exato_1 PORT MAP(
	A=> C(	346	),
	B=> E(	215	),
	Cin=> Carry( 	281	),
	Cout=> Carry( 	282	),
	S=> E(	277	));
			
 U283	: Somador_Exato_1 PORT MAP(
	A=> C(	347	),
	B=> E(	216	),
	Cin=> Carry( 	282	),
	Cout=> Carry( 	283	),
	S=> E(	278	));
			
 U284	: Somador_Exato_1 PORT MAP(
	A=> C(	348	),
	B=> E(	217	),
	Cin=> Carry( 	283	),
	Cout=> Carry( 	284	),
	S=> E(	279	));
			
 U285	: Somador_Exato_1 PORT MAP(
	A=> C(	349	),
	B=> E(	218	),
	Cin=> Carry( 	284	),
	Cout=> Carry( 	285	),
	S=> E(	280	));
			
 U286	: Somador_Exato_1 PORT MAP(
	A=> C(	350	),
	B=> E(	219	),
	Cin=> Carry( 	285	),
	Cout=> Carry( 	286	),
	S=> E(	281	));
			
 U287	: Somador_Exato_1 PORT MAP(
	A=> C(	351	),
	B=> E(	220	),
	Cin=> Carry( 	286	),
	Cout=> Carry( 	287	),
	S=> E(	282	));
			
 U288	: Somador_Exato_1 PORT MAP(
	A=> C(	352	),
	B=> E(	221	),
	Cin=> Carry( 	287	),
	Cout=> Carry( 	288	),
	S=> E(	283	));
			
 U289	: Somador_Exato_1 PORT MAP(
	A=> C(	353	),
	B=> E(	222	),
	Cin=> Carry( 	288	),
	Cout=> Carry( 	289	),
	S=> E(	284	));
			
 U290	: Somador_Exato_1 PORT MAP(
	A=> C(	354	),
	B=> E(	223	),
	Cin=> Carry( 	289	),
	Cout=> Carry( 	290	),
	S=> E(	285	));
			
 U291	: Somador_Exato_1 PORT MAP(
	A=> C(	355	),
	B=> E(	224	),
	Cin=> Carry( 	290	),
	Cout=> Carry( 	291	),
	S=> E(	286	));
			
 U292	: Somador_Exato_1 PORT MAP(
	A=> C(	356	),
	B=> E(	225	),
	Cin=> Carry( 	291	),
	Cout=> Carry( 	292	),
	S=> E(	287	));
			
 U293	: Somador_Exato_1 PORT MAP(
	A=> C(	357	),
	B=> E(	226	),
	Cin=> Carry( 	292	),
	Cout=> Carry( 	293	),
	S=> E(	288	));
			
 U294	: Somador_Exato_1 PORT MAP(
	A=> C(	358	),
	B=> E(	227	),
	Cin=> Carry( 	293	),
	Cout=> Carry( 	294	),
	S=> E(	289	));
			
 U295	: Somador_Exato_1 PORT MAP(
	A=> C(	359	),
	B=> E(	228	),
	Cin=> Carry( 	294	),
	Cout=> Carry( 	295	),
	S=> E(	290	));
			
 U296	: Somador_Exato_1 PORT MAP(
	A=> C(	360	),
	B=> E(	229	),
	Cin=> Carry( 	295	),
	Cout=> Carry( 	296	),
	S=> E(	291	));
			
 U297	: Somador_Exato_1 PORT MAP(
	A=> C(	361	),
	B=> E(	230	),
	Cin=> Carry( 	296	),
	Cout=> Carry( 	297	),
	S=> E(	292	));
			
 U298	: Somador_Exato_1 PORT MAP(
	A=> C(	362	),
	B=> E(	231	),
	Cin=> Carry( 	297	),
	Cout=> Carry( 	298	),
	S=> E(	293	));
			
 U299	: Somador_Exato_1 PORT MAP(
	A=> C(	363	),
	B=> E(	232	),
	Cin=> Carry( 	298	),
	Cout=> Carry( 	299	),
	S=> E(	294	));
			
 U300	: Somador_Exato_1 PORT MAP(
	A=> C(	364	),
	B=> E(	233	),
	Cin=> Carry( 	299	),
	Cout=> Carry( 	300	),
	S=> E(	295	));
			
 U301	: Somador_Exato_1 PORT MAP(
	A=> C(	365	),
	B=> E(	234	),
	Cin=> Carry( 	300	),
	Cout=> Carry( 	301	),
	S=> E(	296	));
			
 U302	: Somador_Exato_1 PORT MAP(
	A=> C(	366	),
	B=> E(	235	),
	Cin=> Carry( 	301	),
	Cout=> Carry( 	302	),
	S=> E(	297	));
			
 U303	: Somador_Exato_1 PORT MAP(
	A=> C(	367	),
	B=> E(	236	),
	Cin=> Carry( 	302	),
	Cout=> Carry( 	303	),
	S=> E(	298	));
			
 U304	: Somador_Exato_1 PORT MAP(
	A=> C(	368	),
	B=> E(	237	),
	Cin=> Carry( 	303	),
	Cout=> Carry( 	304	),
	S=> E(	299	));
			
 U305	: Somador_Exato_1 PORT MAP(
	A=> C(	369	),
	B=> E(	238	),
	Cin=> Carry( 	304	),
	Cout=> Carry( 	305	),
	S=> E(	300	));
			
 U306	: Somador_Exato_1 PORT MAP(
	A=> C(	370	),
	B=> E(	239	),
	Cin=> Carry( 	305	),
	Cout=> Carry( 	306	),
	S=> E(	301	));
			
 U307	: Somador_Exato_1 PORT MAP(
	A=> C(	371	),
	B=> E(	240	),
	Cin=> Carry( 	306	),
	Cout=> Carry( 	307	),
	S=> E(	302	));
			
 U308	: Somador_Exato_1 PORT MAP(
	A=> C(	372	),
	B=> E(	241	),
	Cin=> Carry( 	307	),
	Cout=> Carry( 	308	),
	S=> E(	303	));
			
 U309	: Somador_Exato_1 PORT MAP(
	A=> C(	373	),
	B=> E(	242	),
	Cin=> Carry( 	308	),
	Cout=> Carry( 	309	),
	S=> E(	304	));
			
 U310	: Somador_Exato_1 PORT MAP(
	A=> C(374),
	B=> E(243),
	Cin=> Carry(309),
	Cout=> Carry(310),
	S=> E(305));
			
 U311	: Somador_Exato_1 PORT MAP(
	A=> C(	375	),
	B=> E(	244	),
	Cin=> Carry( 	310	),
	Cout=> Carry( 	311	),
	S=> E(	306	));
			
 U312	: Somador_Exato_1 PORT MAP(
	A=> C(	376	),
	B=> E(	245	),
	Cin=> Carry( 	311	),
	Cout=> Carry( 	312	),
	S=> E(	307	));
			
 U313	: Somador_Exato_1 PORT MAP(
	A=> C(	377	),
	B=> E(	246	),
	Cin=> Carry( 	312	),
	Cout=> Carry( 	313	),
	S=> E(	308	));
			
 U314	: Somador_Exato_1 PORT MAP(
	A=> C(	378	),
	B=> E(	247	),
	Cin=> Carry( 	313	),
	Cout=> Carry( 	314	),
	S=> E(	309	));
			
 U315	: Somador_Exato_1 PORT MAP(
	A=> C(	379	),
	B=> E(	248	),
	Cin=> Carry( 	314	),
	Cout=> Carry( 	315	),
	S=> E(	310	));
			
 U316	: Somador_Exato_1 PORT MAP(
	A=> C(	380	),
	B=> E(	249	),
	Cin=> Carry( 	315	),
	Cout=> Carry( 	316	),
	S=> E(	311	));
			
 U317	: Somador_Exato_1 PORT MAP(
	A=> C(	381	),
	B=> E(	250	),
	Cin=> Carry( 	316	),
	Cout=> Carry( 	317	),
	S=> E(	312	));
			
 U318	: Somador_Exato_1 PORT MAP(
	A=> C(	382	),
	B=> E(	251	),
	Cin=> Carry( 	317	),
	Cout=> Carry( 	318	),
	S=> E(	313	));
			
 U319	: Somador_Exato_1 PORT MAP(
	A => C(383),
	B => Carry(255),
	Cin => Carry(318),
	Cout => Carry(319),
	S => E(314));
---6

			
 U320	: Somador_Exato_1 PORT MAP(
	A=> C(	384	),
	B=> E(	252	),
	Cin=> '0'	,
	Cout=> Carry( 	320	),
	S=> R(	6	));
			
 U321	: Somador_Exato_1 PORT MAP(
	A=> C(	385	),
	B=> E(	253	),
	Cin=> Carry( 	320	),
	Cout=> Carry( 	321	),
	S=> E(	315	));
			
 U322	: Somador_Exato_1 PORT MAP(
	A=> C(	386	),
	B=> E(	254	),
	Cin=> Carry( 	321	),
	Cout=> Carry( 	322	),
	S=> E(	316	));
			
 U323	: Somador_Exato_1 PORT MAP(
	A=> C(	387	),
	B=> E(	255	),
	Cin=> Carry( 	322	),
	Cout=> Carry( 	323	),
	S=> E(	317	));
			
 U324	: Somador_Exato_1 PORT MAP(
	A=> C(	388	),
	B=> E(	256	),
	Cin=> Carry( 	323	),
	Cout=> Carry( 	324	),
	S=> E(	318	));
 			
 U325	: Somador_Exato_1 PORT MAP(
	A=> C(	389	),
	B=> E(	257	),
	Cin=> Carry( 	324	),
	Cout=> Carry( 	325	),
	S=> E(	319	));
			
 U326	: Somador_Exato_1 PORT MAP(
	A=> C(	390	),
	B=> E(	258	),
	Cin=> Carry( 	325	),
	Cout=> Carry( 	326	),
	S=> E(	320	));
			
 U327	: Somador_Exato_1 PORT MAP(
	A=> C(	391	),
	B=> E(	259	),
	Cin=> Carry( 	326	),
	Cout=> Carry( 	327	),
	S=> E(	321	));
			
 U328	: Somador_Exato_1 PORT MAP(
	A=> C(	392	),
	B=> E(	260	),
	Cin=> Carry( 	327	),
	Cout=> Carry( 	328	),
	S=> E(	322	));
			
 U329	: Somador_Exato_1 PORT MAP(
	A=> C(	393	),
	B=> E(	261	),
	Cin=> Carry( 	328	),
	Cout=> Carry( 	329	),
	S=> E(	323	));
			
 U330	: Somador_Exato_1 PORT MAP(
	A=> C(	394	),
	B=> E(	262	),
	Cin=> Carry( 	329	),
	Cout=> Carry( 	330	),
	S=> E(	324	));
			
 U331	: Somador_Exato_1 PORT MAP(
	A=> C(	395	),
	B=> E(	263	),
	Cin=> Carry( 	330	),
	Cout=> Carry( 	331	),
	S=> E(	325	));
			
 U332	: Somador_Exato_1 PORT MAP(
	A=> C(	396	),
	B=> E(	264	),
	Cin=> Carry( 	331	),
	Cout=> Carry( 	332	),
	S=> E(	326	));
			
 U333	: Somador_Exato_1 PORT MAP(
	A=> C(	397	),
	B=> E(	265	),
	Cin=> Carry( 	332	),
	Cout=> Carry( 	333	),
	S=> E(	327	));
			
 U334	: Somador_Exato_1 PORT MAP(
	A=> C(	398	),
	B=> E(	266	),
	Cin=> Carry( 	333	),
	Cout=> Carry( 	334	),
	S=> E(	328	));
			
 U335	: Somador_Exato_1 PORT MAP(
	A=> C(	399	),
	B=> E(	267	),
	Cin=> Carry( 	334	),
	Cout=> Carry( 	335	),
	S=> E(	329	));
			
 U336	: Somador_Exato_1 PORT MAP(
	A=> C(	400	),
	B=> E(	268	),
	Cin=> Carry( 	335	),
	Cout=> Carry( 	336	),
	S=> E(	330	));
			
 U337	: Somador_Exato_1 PORT MAP(
	A=> C(	401	),
	B=> E(	269	),
	Cin=> Carry( 	336	),
	Cout=> Carry( 	337	),
	S=> E(	331	));
			
 U338	: Somador_Exato_1 PORT MAP(
	A=> C(	402	),
	B=> E(	270	),
	Cin=> Carry( 	337	),
	Cout=> Carry( 	338	),
	S=> E(	332	));
			
 U339	: Somador_Exato_1 PORT MAP(
	A=> C(	403	),
	B=> E(	271	),
	Cin=> Carry( 	338	),
	Cout=> Carry( 	339	),
	S=> E(	333	));
			
 U340	: Somador_Exato_1 PORT MAP(
	A=> C(	404	),
	B=> E(	272	),
	Cin=> Carry( 	339	),
	Cout=> Carry( 	340	),
	S=> E(	334	));
			
 U341	: Somador_Exato_1 PORT MAP(
	A=> C(	405	),
	B=> E(	273	),
	Cin=> Carry( 	340	),
	Cout=> Carry( 	341	),
	S=> E(	335	));
			
 U342	: Somador_Exato_1 PORT MAP(
	A=> C(	406	),
	B=> E(	274	),
	Cin=> Carry( 	341	),
	Cout=> Carry( 	342	),
	S=> E(	336	));
			
 U343	: Somador_Exato_1 PORT MAP(
	A=> C(	407	),
	B=> E(	275	),
	Cin=> Carry( 	342	),
	Cout=> Carry( 	343	),
	S=> E(	337	));
			
 U344	: Somador_Exato_1 PORT MAP(
	A=> C(	408	),
	B=> E(	276	),
	Cin=> Carry( 	343	),
	Cout=> Carry( 	344	),
	S=> E(	338	));
			
 U345	: Somador_Exato_1 PORT MAP(
	A=> C(	409	),
	B=> E(	277	),
	Cin=> Carry( 	344	),
	Cout=> Carry( 	345	),
	S=> E(	339	));
			
 U346	: Somador_Exato_1 PORT MAP(
	A=> C(	410	),
	B=> E(	278	),
	Cin=> Carry( 	345	),
	Cout=> Carry( 	346	),
	S=> E(	340	));
			
 U347	: Somador_Exato_1 PORT MAP(
	A=> C(	411	),
	B=> E(	279	),
	Cin=> Carry( 	346	),
	Cout=> Carry( 	347	),
	S=> E(	341	));
			
 U348	: Somador_Exato_1 PORT MAP(
	A=> C(	412	),
	B=> E(	280	),
	Cin=> Carry( 	347	),
	Cout=> Carry( 	348	),
	S=> E(	342	));
			
 U349	: Somador_Exato_1 PORT MAP(
	A=> C(	413	),
	B=> E(	281	),
	Cin=> Carry( 	348	),
	Cout=> Carry( 	349	),
	S=> E(	343	));
			
 U350	: Somador_Exato_1 PORT MAP(
	A=> C(	414	),
	B=> E(	282	),
	Cin=> Carry( 	349	),
	Cout=> Carry( 	350	),
	S=> E(	344	));
			
 U351	: Somador_Exato_1 PORT MAP(
	A=> C(	415	),
	B=> E(	283	),
	Cin=> Carry( 	350	),
	Cout=> Carry( 	351	),
	S=> E(	345	));
			
 U352	: Somador_Exato_1 PORT MAP(
	A=> C(	416	),
	B=> E(	284	),
	Cin=> Carry( 	351	),
	Cout=> Carry( 	352	),
	S=> E(	346	));
			
 U353	: Somador_Exato_1 PORT MAP(
	A=> C(	417	),
	B=> E(	285	),
	Cin=> Carry( 	352	),
	Cout=> Carry( 	353	),
	S=> E(	347	));
			
 U354	: Somador_Exato_1 PORT MAP(
	A=> C(	418	),
	B=> E(	286	),
	Cin=> Carry( 	353	),
	Cout=> Carry( 	354	),
	S=> E(	348	));
			
 U355	: Somador_Exato_1 PORT MAP(
	A=> C(	419	),
	B=> E(	287	),
	Cin=> Carry( 	354	),
	Cout=> Carry( 	355	),
	S=> E(	349	));
			
 U356	: Somador_Exato_1 PORT MAP(
	A=> C(	420	),
	B=> E(	288	),
	Cin=> Carry( 	355	),
	Cout=> Carry( 	356	),
	S=> E(	350	));
			
 U357	: Somador_Exato_1 PORT MAP(
	A=> C(	421	),
	B=> E(	289	),
	Cin=> Carry( 	356	),
	Cout=> Carry( 	357	),
	S=> E(	351	));
			
 U358	: Somador_Exato_1 PORT MAP(
	A=> C(	422	),
	B=> E(	290	),
	Cin=> Carry( 	357	),
	Cout=> Carry( 	358	),
	S=> E(	352	));
			
 U359	: Somador_Exato_1 PORT MAP(
	A=> C(	423	),
	B=> E(	291	),
	Cin=> Carry( 	358	),
	Cout=> Carry( 	359	),
	S=> E(	353	));
			
 U360	: Somador_Exato_1 PORT MAP(
	A=> C(	424	),
	B=> E(	292	),
	Cin=> Carry( 	359	),
	Cout=> Carry( 	360	),
	S=> E(	354	));
			
 U361	: Somador_Exato_1 PORT MAP(
	A=> C(	425	),
	B=> E(	293	),
	Cin=> Carry( 	360	),
	Cout=> Carry( 	361	),
	S=> E(	355	));
			
 U362	: Somador_Exato_1 PORT MAP(
	A=> C(	426	),
	B=> E(	294	),
	Cin=> Carry( 	361	),
	Cout=> Carry( 	362	),
	S=> E(	356	));
			
 U363	: Somador_Exato_1 PORT MAP(
	A=> C(	427	),
	B=> E(	295	),
	Cin=> Carry( 	362	),
	Cout=> Carry( 	363	),
	S=> E(	357	));
			
 U364	: Somador_Exato_1 PORT MAP(
	A=> C(	428	),
	B=> E(	296	),
	Cin=> Carry( 	363	),
	Cout=> Carry( 	364	),
	S=> E(	358	));
			
 U365	: Somador_Exato_1 PORT MAP(
	A=> C(	429	),
	B=> E(	297	),
	Cin=> Carry( 	364	),
	Cout=> Carry( 	365	),
	S=> E(	359	));
			
 U366	: Somador_Exato_1 PORT MAP(
	A=> C(	430	),
	B=> E(	298	),
	Cin=> Carry( 	365	),
	Cout=> Carry( 	366	),
	S=> E(	360	));
			
 U367	: Somador_Exato_1 PORT MAP(
	A=> C(	431	),
	B=> E(	299	),
	Cin=> Carry( 	366	),
	Cout=> Carry( 	367	),
	S=> E(	361	));
			
 U368	: Somador_Exato_1 PORT MAP(
	A=> C(	432	),
	B=> E(	300	),
	Cin=> Carry( 	367	),
	Cout=> Carry( 	368	),
	S=> E(	362	));
			
 U369	: Somador_Exato_1 PORT MAP(
	A=> C(	433	),
	B=> E(	301	),
	Cin=> Carry( 	368	),
	Cout=> Carry( 	369	),
	S=> E(	363	));
			
 U370	: Somador_Exato_1 PORT MAP(
	A=> C(	434	),
	B=> E(	302	),
	Cin=> Carry( 	369	),
	Cout=> Carry( 	370	),
	S=> E(	364	));
			
 U371	: Somador_Exato_1 PORT MAP(
	A=> C(	435	),
	B=> E(	303	),
	Cin=> Carry( 	370	),
	Cout=> Carry( 	371	),
	S=> E(	365	));
			
 U372	: Somador_Exato_1 PORT MAP(
	A=> C(	436	),
	B=> E(	304	),
	Cin=> Carry( 	371	),
	Cout=> Carry( 	372	),
	S=> E(	366	));
			
 U373	: Somador_Exato_1 PORT MAP(
	A=> C(	437	),
	B=> E(	305	),
	Cin=> Carry( 	372	),
	Cout=> Carry( 	373	),
	S=> E(	367	));
			
 U374	: Somador_Exato_1 PORT MAP(
	A=> C(	438	),
	B=> E(	306	),
	Cin=> Carry( 	373	),
	Cout=> Carry( 	374	),
	S=> E(	368	));
			
 U375	: Somador_Exato_1 PORT MAP(
	A=> C(	439	),
	B=> E(	307	),
	Cin=> Carry( 	374	),
	Cout=> Carry( 	375	),
	S=> E(	369	));
			
 U376	: Somador_Exato_1 PORT MAP(
	A=> C(	440	),
	B=> E(	308	),
	Cin=> Carry( 	375	),
	Cout=> Carry( 	376	),
	S=> E(	370	));
			
 U377	: Somador_Exato_1 PORT MAP(
	A=> C(	441	),
	B=> E(	309	),
	Cin=> Carry( 	376	),
	Cout=> Carry( 	377	),
	S=> E(	371	));
			
 U378	: Somador_Exato_1 PORT MAP(
	A=> C(	442	),
	B=> E(	310	),
	Cin=> Carry( 	377	),
	Cout=> Carry( 	378	),
	S=> E(	372	));
			
 U379	: Somador_Exato_1 PORT MAP(
	A=> C(	443	),
	B=> E(	311	),
	Cin=> Carry( 	378	),
	Cout=> Carry( 	379	),
	S=> E(	373	));
			
 U380	: Somador_Exato_1 PORT MAP(
	A=> C(	444	),
	B=> E(	312	),
	Cin=> Carry( 	379	),
	Cout=> Carry( 	380	),
	S=> E(	374	));
			
 U381	: Somador_Exato_1 PORT MAP(
	A=> C(	445	),
	B=> E(	313	),
	Cin=> Carry( 	380	),
	Cout=> Carry( 	381	),
	S=> E(	375	));
			
 U382	: Somador_Exato_1 PORT MAP(
	A=> C(	446	),
	B=> E(	314	),
	Cin=> Carry( 	381	),
	Cout=> Carry( 	382	),
	S=> E(	376	));
			
 U383	: Somador_Exato_1 PORT MAP(
	A=> C(	447	),
	B=> Carry(	319	),
	Cin=> Carry( 	382	),
	Cout=> Carry( 	383	),
	S=> E(	377	));

----

			
 U384	: Somador_Exato_1 PORT MAP(
	A=> C(	448	),
	B=> E(	315	),
	Cin=> '0'	,
	Cout=> Carry( 	384	),
	S=> R(	7	));
			
 U385	: Somador_Exato_1 PORT MAP(
	A=> C(	449	),
	B=> E(	316	),
	Cin=> Carry( 	384	),
	Cout=> Carry( 	385	),
	S=> E(	378	));
			
 U386	: Somador_Exato_1 PORT MAP(
	A=> C(	450	),
	B=> E(	317	),
	Cin=> Carry( 	385	),
	Cout=> Carry( 	386	),
	S=> E(	379	));
			
 U387	: Somador_Exato_1 PORT MAP(
	A=> C(	451	),
	B=> E(	318	),
	Cin=> Carry( 	386	),
	Cout=> Carry( 	387	),
	S=> E(	380	));
			
 U388	: Somador_Exato_1 PORT MAP(
	A=> C(	452	),
	B=> E(	319	),
	Cin=> Carry( 	387	),
	Cout=> Carry( 	388	),
	S=> E(	381	));
			
 U389	: Somador_Exato_1 PORT MAP(
	A=> C(	453	),
	B=> E(	320	),
	Cin=> Carry( 	388	),
	Cout=> Carry( 	389	),
	S=> E(	382	));
			
 U390	: Somador_Exato_1 PORT MAP(
	A=> C(	454	),
	B=> E(	321	),
	Cin=> Carry( 	389	),
	Cout=> Carry( 	390	),
	S=> E(	383	));
			
 U391	: Somador_Exato_1 PORT MAP(
	A=> C(	455	),
	B=> E(	322	),
	Cin=> Carry( 	390	),
	Cout=> Carry( 	391	),
	S=> E(	384	));
			
 U392	: Somador_Exato_1 PORT MAP(
	A=> C(	456	),
	B=> E(	323	),
	Cin=> Carry( 	391	),
	Cout=> Carry( 	392	),
	S=> E(	385	));
			
 U393	: Somador_Exato_1 PORT MAP(
	A=> C(	457	),
	B=> E(	324	),
	Cin=> Carry( 	392	),
	Cout=> Carry( 	393	),
	S=> E(	386	));
			
 U394	: Somador_Exato_1 PORT MAP(
	A=> C(	458	),
	B=> E(	325	),
	Cin=> Carry( 	393	),
	Cout=> Carry( 	394	),
	S=> E(	387	));
			
 U395	: Somador_Exato_1 PORT MAP(
	A=> C(	459	),
	B=> E(	326	),
	Cin=> Carry( 	394	),
	Cout=> Carry( 	395	),
	S=> E(	388	));
			
 U396	: Somador_Exato_1 PORT MAP(
	A=> C(	460	),
	B=> E(	327	),
	Cin=> Carry( 	395	),
	Cout=> Carry( 	396	),
	S=> E(	389	));
			
 U397	: Somador_Exato_1 PORT MAP(
	A=> C(	461	),
	B=> E(	328	),
	Cin=> Carry( 	396	),
	Cout=> Carry( 	397	),
	S=> E(	390	));
			
 U398	: Somador_Exato_1 PORT MAP(
	A=> C(	462	),
	B=> E(	329	),
	Cin=> Carry( 	397	),
	Cout=> Carry( 	398	),
	S=> E(	391	));
			
 U399	: Somador_Exato_1 PORT MAP(
	A=> C(	463	),
	B=> E(	330	),
	Cin=> Carry( 	398	),
	Cout=> Carry( 	399	),
	S=> E(	392	));
			
 U400	: Somador_Exato_1 PORT MAP(
	A=> C(	464	),
	B=> E(	331	),
	Cin=> Carry( 	399	),
	Cout=> Carry( 	400	),
	S=> E(	393	));
			
 U401	: Somador_Exato_1 PORT MAP(
	A=> C(	465	),
	B=> E(	332	),
	Cin=> Carry( 	400	),
	Cout=> Carry( 	401	),
	S=> E(	394	));
			
 U402	: Somador_Exato_1 PORT MAP(
	A=> C(	466	),
	B=> E(	333	),
	Cin=> Carry( 	401	),
	Cout=> Carry( 	402	),
	S=> E(	395	));
			
 U403	: Somador_Exato_1 PORT MAP(
	A=> C(	467	),
	B=> E(	334	),
	Cin=> Carry( 	402	),
	Cout=> Carry( 	403	),
	S=> E(	396	));
			
 U404	: Somador_Exato_1 PORT MAP(
	A=> C(	468	),
	B=> E(	335	),
	Cin=> Carry( 	403	),
	Cout=> Carry( 	404	),
	S=> E(	397	));
			
 U405	: Somador_Exato_1 PORT MAP(
	A=> C(	469	),
	B=> E(	336	),
	Cin=> Carry( 	404	),
	Cout=> Carry( 	405	),
	S=> E(	398	));
			
 U406	: Somador_Exato_1 PORT MAP(
	A=> C(	470	),
	B=> E(	337	),
	Cin=> Carry( 	405	),
	Cout=> Carry( 	406	),
	S=> E(	399	));
			
 U407	: Somador_Exato_1 PORT MAP(
	A=> C(	471	),
	B=> E(	338	),
	Cin=> Carry( 	406	),
	Cout=> Carry( 	407	),
	S=> E(	400	));
			
 U408	: Somador_Exato_1 PORT MAP(
	A=> C(	472	),
	B=> E(	339	),
	Cin=> Carry( 	407	),
	Cout=> Carry( 	408	),
	S=> E(	401	));
			
 U409	: Somador_Exato_1 PORT MAP(
	A=> C(	473	),
	B=> E(	340	),
	Cin=> Carry( 	408	),
	Cout=> Carry( 	409	),
	S=> E(	402	));
			
 U410	: Somador_Exato_1 PORT MAP(
	A=> C(	474	),
	B=> E(	341	),
	Cin=> Carry( 	409	),
	Cout=> Carry( 	410	),
	S=> E(	403	));
			
 U411	: Somador_Exato_1 PORT MAP(
	A=> C(	475	),
	B=> E(	342	),
	Cin=> Carry( 	410	),
	Cout=> Carry( 	411	),
	S=> E(	404	));
			
 U412	: Somador_Exato_1 PORT MAP(
	A=> C(	476	),
	B=> E(	343	),
	Cin=> Carry( 	411	),
	Cout=> Carry( 	412	),
	S=> E(	405	));
			
 U413	: Somador_Exato_1 PORT MAP(
	A=> C(	477	),
	B=> E(	344	),
	Cin=> Carry( 	412	),
	Cout=> Carry( 	413	),
	S=> E(	406	));
			
 U414	: Somador_Exato_1 PORT MAP(
	A=> C(	478	),
	B=> E(	345	),
	Cin=> Carry( 	413	),
	Cout=> Carry( 	414	),
	S=> E(	407	));
			
 U415	: Somador_Exato_1 PORT MAP(
	A=> C(	479	),
	B=> E(	346	),
	Cin=> Carry( 	414	),
	Cout=> Carry( 	415	),
	S=> E(	408	));
			
 U416	: Somador_Exato_1 PORT MAP(
	A=> C(	480	),
	B=> E(	347	),
	Cin=> Carry( 	415	),
	Cout=> Carry( 	416	),
	S=> E(	409	));
			
 U417	: Somador_Exato_1 PORT MAP(
	A=> C(	481	),
	B=> E(	348	),
	Cin=> Carry( 	416	),
	Cout=> Carry( 	417	),
	S=> E(	410	));
			
 U418	: Somador_Exato_1 PORT MAP(
	A=> C(	482	),
	B=> E(	349	),
	Cin=> Carry( 	417	),
	Cout=> Carry( 	418	),
	S=> E(	411	));
			
 U419	: Somador_Exato_1 PORT MAP(
	A=> C(	483	),
	B=> E(	350	),
	Cin=> Carry( 	418	),
	Cout=> Carry( 	419	),
	S=> E(	412	));
			
 U420	: Somador_Exato_1 PORT MAP(
	A=> C(	484	),
	B=> E(	351	),
	Cin=> Carry( 	419	),
	Cout=> Carry( 	420	),
	S=> E(	413	));
			
 U421	: Somador_Exato_1 PORT MAP(
	A=> C(	485	),
	B=> E(	352	),
	Cin=> Carry( 	420	),
	Cout=> Carry( 	421	),
	S=> E(	414	));
			
 U422	: Somador_Exato_1 PORT MAP(
	A=> C(	486	),
	B=> E(	353	),
	Cin=> Carry( 	421	),
	Cout=> Carry( 	422	),
	S=> E(	415	));
			
 U423	: Somador_Exato_1 PORT MAP(
	A=> C(	487	),
	B=> E(	354	),
	Cin=> Carry( 	422	),
	Cout=> Carry( 	423	),
	S=> E(	416	));
			
 U424	: Somador_Exato_1 PORT MAP(
	A=> C(	488	),
	B=> E(	355	),
	Cin=> Carry( 	423	),
	Cout=> Carry( 	424	),
	S=> E(	417	));
			
 U425	: Somador_Exato_1 PORT MAP(
	A=> C(	489	),
	B=> E(	356	),
	Cin=> Carry( 	424	),
	Cout=> Carry( 	425	),
	S=> E(	418	));
			
 U426	: Somador_Exato_1 PORT MAP(
	A=> C(	490	),
	B=> E(	357	),
	Cin=> Carry( 	425	),
	Cout=> Carry( 	426	),
	S=> E(	419	));
			
 U427	: Somador_Exato_1 PORT MAP(
	A=> C(	491	),
	B=> E(	358	),
	Cin=> Carry( 	426	),
	Cout=> Carry( 	427	),
	S=> E(	420	));
			
 U428	: Somador_Exato_1 PORT MAP(
	A=> C(	492	),
	B=> E(	359	),
	Cin=> Carry( 	427	),
	Cout=> Carry( 	428	),
	S=> E(	421	));
			
 U429	: Somador_Exato_1 PORT MAP(
	A=> C(	493	),
	B=> E(	360	),
	Cin=> Carry( 	428	),
	Cout=> Carry( 	429	),
	S=> E(	422	));
			
 U430	: Somador_Exato_1 PORT MAP(
	A=> C(	494	),
	B=> E(	361	),
	Cin=> Carry( 	429	),
	Cout=> Carry( 	430	),
	S=> E(	423	));
			
 U431	: Somador_Exato_1 PORT MAP(
	A=> C(	495	),
	B=> E(	362	),
	Cin=> Carry( 	430	),
	Cout=> Carry( 	431	),
	S=> E(	424	));
			
 U432	: Somador_Exato_1 PORT MAP(
	A=> C(	496	),
	B=> E(	363	),
	Cin=> Carry( 	431	),
	Cout=> Carry( 	432	),
	S=> E(	425	));
			
 U433	: Somador_Exato_1 PORT MAP(
	A=> C(	497	),
	B=> E(	364	),
	Cin=> Carry( 	432	),
	Cout=> Carry( 	433	),
	S=> E(	426	));
			
 U434	: Somador_Exato_1 PORT MAP(
	A=> C(	498	),
	B=> E(	365	),
	Cin=> Carry( 	433	),
	Cout=> Carry( 	434	),
	S=> E(	427	));
			
 U435	: Somador_Exato_1 PORT MAP(
	A=> C(	499	),
	B=> E(	366	),
	Cin=> Carry( 	434	),
	Cout=> Carry( 	435	),
	S=> E(	428	));
			
 U436	: Somador_Exato_1 PORT MAP(
	A=> C(	500	),
	B=> E(	367	),
	Cin=> Carry( 	435	),
	Cout=> Carry( 	436	),
	S=> E(	429	));
			
 U437	: Somador_Exato_1 PORT MAP(
	A=> C(	501	),
	B=> E(	368	),
	Cin=> Carry( 	436	),
	Cout=> Carry( 	437	),
	S=> E(	430	));
			
 U438	: Somador_Exato_1 PORT MAP(
	A=> C(	502	),
	B=> E(	369	),
	Cin=> Carry( 	437	),
	Cout=> Carry( 	438	),
	S=> E(	431	));
			
 U439	: Somador_Exato_1 PORT MAP(
	A=> C(	503	),
	B=> E(	370	),
	Cin=> Carry( 	438	),
	Cout=> Carry( 	439	),
	S=> E(	432	));
			
 U440	: Somador_Exato_1 PORT MAP(
	A=> C(	504	),
	B=> E(	371	),
	Cin=> Carry( 	439	),
	Cout=> Carry( 	440	),
	S=> E(	433	));
			
 U441	: Somador_Exato_1 PORT MAP(
	A=> C(	505	),
	B=> E(	372	),
	Cin=> Carry( 	440	),
	Cout=> Carry( 	441	),
	S=> E(	434	));
			
 U442	: Somador_Exato_1 PORT MAP(
	A=> C(	506	),
	B=> E(	373	),
	Cin=> Carry( 	441	),
	Cout=> Carry( 	442	),
	S=> E(	435	));
			
 U443	: Somador_Exato_1 PORT MAP(
	A=> C(	507	),
	B=> E(	374	),
	Cin=> Carry( 	442	),
	Cout=> Carry( 	443	),
	S=> E(	436	));
			
 U444	: Somador_Exato_1 PORT MAP(
	A=> C(	508	),
	B=> E(	375	),
	Cin=> Carry( 	443	),
	Cout=> Carry( 	444	),
	S=> E(	437	));
			
 U445	: Somador_Exato_1 PORT MAP(
	A=> C(	509	),
	B=> E(	376	),
	Cin=> Carry( 	444	),
	Cout=> Carry( 	445	),
	S=> E(	438	));
			
 U446	: Somador_Exato_1 PORT MAP(
	A=> C(	510	),
	B=> E(	377	),
	Cin=> Carry( 	445	),
	Cout=> Carry( 	446	),
	S=> E(	439	));
			
 U447	: Somador_Exato_1 PORT MAP(
	A=> C(	511	),
	B=> Carry(	383	),
	Cin=> Carry( 	446	),
	Cout=> Carry( 	447	),
	S=> E(	440	));
---
			
 U448	: Somador_Exato_1 PORT MAP(
	A=> C(	512	),
	B=> E(	378	),
	Cin=> '0'	,
	Cout=> Carry( 	448	),
	S=> R(	8	));
			
 U449	: Somador_Exato_1 PORT MAP(
	A=> C(	513	),
	B=> E(	379	),
	Cin=> Carry( 	448	),
	Cout=> Carry( 	449	),
	S=> E(	441	));
			
 U450	: Somador_Exato_1 PORT MAP(
	A=> C(	514	),
	B=> E(	380	),
	Cin=> Carry( 	449	),
	Cout=> Carry( 	450	),
	S=> E(	442	));
			
 U451	: Somador_Exato_1 PORT MAP(
	A=> C(	515	),
	B=> E(	381	),
	Cin=> Carry( 	450	),
	Cout=> Carry( 	451	),
	S=> E(	443	));
			
 U452	: Somador_Exato_1 PORT MAP(
	A=> C(	516	),
	B=> E(	382	),
	Cin=> Carry( 	451	),
	Cout=> Carry( 	452	),
	S=> E(	444	));
			
 U453	: Somador_Exato_1 PORT MAP(
	A=> C(	517	),
	B=> E(	383	),
	Cin=> Carry( 	452	),
	Cout=> Carry( 	453	),
	S=> E(	445	));
			
 U454	: Somador_Exato_1 PORT MAP(
	A=> C(	518	),
	B=> E(	384	),
	Cin=> Carry( 	453	),
	Cout=> Carry( 	454	),
	S=> E(	446	));
			
 U455	: Somador_Exato_1 PORT MAP(
	A=> C(	519	),
	B=> E(	385	),
	Cin=> Carry( 	454	),
	Cout=> Carry( 	455	),
	S=> E(	447	));
			
 U456	: Somador_Exato_1 PORT MAP(
	A=> C(	520	),
	B=> E(	386	),
	Cin=> Carry( 	455	),
	Cout=> Carry( 	456	),
	S=> E(	448	));
			
 U457	: Somador_Exato_1 PORT MAP(
	A=> C(	521	),
	B=> E(	387	),
	Cin=> Carry( 	456	),
	Cout=> Carry( 	457	),
	S=> E(	449	));
			
 U458	: Somador_Exato_1 PORT MAP(
	A=> C(	522	),
	B=> E(	388	),
	Cin=> Carry( 	457	),
	Cout=> Carry( 	458	),
	S=> E(	450	));
			
 U459	: Somador_Exato_1 PORT MAP(
	A=> C(	523	),
	B=> E(	389	),
	Cin=> Carry( 	458	),
	Cout=> Carry( 	459	),
	S=> E(	451	));
			
 U460	: Somador_Exato_1 PORT MAP(
	A=> C(	524	),
	B=> E(	390	),
	Cin=> Carry( 	459	),
	Cout=> Carry( 	460	),
	S=> E(	452	));
			
 U461	: Somador_Exato_1 PORT MAP(
	A=> C(	525	),
	B=> E(	391	),
	Cin=> Carry( 	460	),
	Cout=> Carry( 	461	),
	S=> E(	453	));
			
 U462	: Somador_Exato_1 PORT MAP(
	A=> C(	526	),
	B=> E(	392	),
	Cin=> Carry( 	461	),
	Cout=> Carry( 	462	),
	S=> E(	454	));
			
 U463	: Somador_Exato_1 PORT MAP(
	A=> C(	527	),
	B=> E(	393	),
	Cin=> Carry( 	462	),
	Cout=> Carry( 	463	),
	S=> E(	455	));
			
 U464	: Somador_Exato_1 PORT MAP(
	A=> C(	528	),
	B=> E(	394	),
	Cin=> Carry( 	463	),
	Cout=> Carry( 	464	),
	S=> E(	456	));
			
 U465	: Somador_Exato_1 PORT MAP(
	A=> C(	529	),
	B=> E(	395	),
	Cin=> Carry( 	464	),
	Cout=> Carry( 	465	),
	S=> E(	457	));
			
 U466	: Somador_Exato_1 PORT MAP(
	A=> C(	530	),
	B=> E(	396	),
	Cin=> Carry( 	465	),
	Cout=> Carry( 	466	),
	S=> E(	458	));
			
 U467	: Somador_Exato_1 PORT MAP(
	A=> C(	531	),
	B=> E(	397	),
	Cin=> Carry( 	466	),
	Cout=> Carry( 	467	),
	S=> E(	459	));
			
U468	: Somador_Exato_1 PORT MAP(
	A=> C(	532	),
	B=> E(	398	),
	Cin=> Carry( 	467	),
	Cout=> Carry( 	468	),
	S=> E(	460	));
			
 U469	: Somador_Exato_1 PORT MAP(
	A=> C(	533	),
	B=> E(	399	),
	Cin=> Carry( 	468	),
	Cout=> Carry( 	469	),
	S=> E(	461	));
			
 U470	: Somador_Exato_1 PORT MAP(
	A=> C(	534	),
	B=> E(	400	),
	Cin=> Carry( 	469	),
	Cout=> Carry( 	470	),
	S=> E(	462	));
			
 U471	: Somador_Exato_1 PORT MAP(
	A=> C(	535	),
	B=> E(	401	),
	Cin=> Carry( 	470	),
	Cout=> Carry( 	471	),
	S=> E(	463	));
			
 U472	: Somador_Exato_1 PORT MAP(
	A=> C(	536	),
	B=> E(	402	),
	Cin=> Carry( 	471	),
	Cout=> Carry( 	472	),
	S=> E(	464	));
			
 U473	: Somador_Exato_1 PORT MAP(
	A=> C(	537	),
	B=> E(	403	),
	Cin=> Carry( 	472	),
	Cout=> Carry( 	473	),
	S=> E(	465	));
			
 U474	: Somador_Exato_1 PORT MAP(
	A=> C(	538	),
	B=> E(	404	),
	Cin=> Carry( 	473	),
	Cout=> Carry( 	474	),
	S=> E(	466	));
			
 U475	: Somador_Exato_1 PORT MAP(
	A=> C(	539	),
	B=> E(	405	),
	Cin=> Carry( 	474	),
	Cout=> Carry( 	475	),
	S=> E(	467	));
			
 U476	: Somador_Exato_1 PORT MAP(
	A=> C(	540	),
	B=> E(	406	),
	Cin=> Carry( 	475	),
	Cout=> Carry( 	476	),
	S=> E(	468	));
			
 U477	: Somador_Exato_1 PORT MAP(
	A=> C(	541	),
	B=> E(	407	),
	Cin=> Carry( 	476	),
	Cout=> Carry( 	477	),
	S=> E(	469	));
			
 U478	: Somador_Exato_1 PORT MAP(
	A=> C(	542	),
	B=> E(	408	),
	Cin=> Carry( 	477	),
	Cout=> Carry( 	478	),
	S=> E(	470	));
			
 U479	: Somador_Exato_1 PORT MAP(
	A=> C(	543	),
	B=> E(	409	),
	Cin=> Carry( 	478	),
	Cout=> Carry( 	479	),
	S=> E(	471	));
			
 U480	: Somador_Exato_1 PORT MAP(
	A=> C(	544	),
	B=> E(	410	),
	Cin=> Carry( 	479	),
	Cout=> Carry( 	480	),
	S=> E(	472	));
			
 U481	: Somador_Exato_1 PORT MAP(
	A=> C(	545	),
	B=> E(	411	),
	Cin=> Carry( 	480	),
	Cout=> Carry( 	481	),
	S=> E(	473	));
			
 U482	: Somador_Exato_1 PORT MAP(
	A=> C(	546	),
	B=> E(	412	),
	Cin=> Carry( 	481	),
	Cout=> Carry( 	482	),
	S=> E(	474	));
			
 U483	: Somador_Exato_1 PORT MAP(
	A=> C(	547	),
	B=> E(	413	),
	Cin=> Carry( 	482	),
	Cout=> Carry( 	483	),
	S=> E(	475	));
			
 U484	: Somador_Exato_1 PORT MAP(
	A=> C(	548	),
	B=> E(	414	),
	Cin=> Carry( 	483	),
	Cout=> Carry( 	484	),
	S=> E(	476	));
			
 U485	: Somador_Exato_1 PORT MAP(
	A=> C(	549	),
	B=> E(	415	),
	Cin=> Carry( 	484	),
	Cout=> Carry( 	485	),
	S=> E(	477	));
			
 U486	: Somador_Exato_1 PORT MAP(
	A=> C(	550	),
	B=> E(	416	),
	Cin=> Carry( 	485	),
	Cout=> Carry( 	486	),
	S=> E(	478	));
			
 U487	: Somador_Exato_1 PORT MAP(
	A=> C(	551	),
	B=> E(	417	),
	Cin=> Carry( 	486	),
	Cout=> Carry( 	487	),
	S=> E(	479	));
			
 U488	: Somador_Exato_1 PORT MAP(
	A=> C(	552	),
	B=> E(	418	),
	Cin=> Carry( 	487	),
	Cout=> Carry( 	488	),
	S=> E(	480	));
			
 U489	: Somador_Exato_1 PORT MAP(
	A=> C(	553	),
	B=> E(	419	),
	Cin=> Carry( 	488	),
	Cout=> Carry( 	489	),
	S=> E(	481	));
			
 U490	: Somador_Exato_1 PORT MAP(
	A=> C(	554	),
	B=> E(	420	),
	Cin=> Carry( 	489	),
	Cout=> Carry( 	490	),
	S=> E(	482	));
			
 U491	: Somador_Exato_1 PORT MAP(
	A=> C(	555	),
	B=> E(	421	),
	Cin=> Carry( 	490	),
	Cout=> Carry( 	491	),
	S=> E(	483	));
			
 U492	: Somador_Exato_1 PORT MAP(
	A=> C(	556	),
	B=> E(	422	),
	Cin=> Carry( 	491	),
	Cout=> Carry( 	492	),
	S=> E(	484	));
			
 U493	: Somador_Exato_1 PORT MAP(
	A=> C(	557	),
	B=> E(	423	),
	Cin=> Carry( 	492	),
	Cout=> Carry( 	493	),
	S=> E(	485	));
			
 U494	: Somador_Exato_1 PORT MAP(
	A=> C(	558	),
	B=> E(	424	),
	Cin=> Carry( 	493	),
	Cout=> Carry( 	494	),
	S=> E(	486	));
			
 U495	: Somador_Exato_1 PORT MAP(
	A=> C(	559	),
	B=> E(	425	),
	Cin=> Carry( 	494	),
	Cout=> Carry( 	495	),
	S=> E(	487	));
			
 U496	: Somador_Exato_1 PORT MAP(
	A=> C(	560	),
	B=> E(	426	),
	Cin=> Carry( 	495	),
	Cout=> Carry( 	496	),
	S=> E(	488	));
			
 U497	: Somador_Exato_1 PORT MAP(
	A=> C(	561	),
	B=> E(	427	),
	Cin=> Carry( 	496	),
	Cout=> Carry( 	497	),
	S=> E(	489	));
			
 U498	: Somador_Exato_1 PORT MAP(
	A=> C(	562	),
	B=> E(	428	),
	Cin=> Carry( 	497	),
	Cout=> Carry( 	498	),
	S=> E(	490	));
			
 U499	: Somador_Exato_1 PORT MAP(
	A=> C(	563	),
	B=> E(	429	),
	Cin=> Carry( 	498	),
	Cout=> Carry( 	499	),
	S=> E(	491	));
			
 U500	: Somador_Exato_1 PORT MAP(
	A=> C(	564	),
	B=> E(	430	),
	Cin=> Carry( 	499	),
	Cout=> Carry( 	500	),
	S=> E(	492	));
			
 U501	: Somador_Exato_1 PORT MAP(
	A=> C(	565	),
	B=> E(	431	),
	Cin=> Carry( 	500	),
	Cout=> Carry( 	501	),
	S=> E(	493	));
			
 U502	: Somador_Exato_1 PORT MAP(
	A=> C(	566	),
	B=> E(	432	),
	Cin=> Carry( 	501	),
	Cout=> Carry( 	502	),
	S=> E(	494	));
			
 U503	: Somador_Exato_1 PORT MAP(
	A=> C(	567	),
	B=> E(	433	),
	Cin=> Carry( 	502	),
	Cout=> Carry( 	503	),
	S=> E(	495	));
			
 U504	: Somador_Exato_1 PORT MAP(
	A=> C(	568	),
	B=> E(	434	),
	Cin=> Carry( 	503	),
	Cout=> Carry( 	504	),
	S=> E(	496	));
			
 U505	: Somador_Exato_1 PORT MAP(
	A=> C(	569	),
	B=> E(	435	),
	Cin=> Carry( 	504	),
	Cout=> Carry( 	505	),
	S=> E(	497	));
			
 U506	: Somador_Exato_1 PORT MAP(
	A=> C(	570	),
	B=> E(	436	),
	Cin=> Carry( 	505	),
	Cout=> Carry( 	506	),
	S=> E(	498	));
			
 U507	: Somador_Exato_1 PORT MAP(
	A=> C(	571	),
	B=> E(	437	),
	Cin=> Carry( 	506	),
	Cout=> Carry( 	507	),
	S=> E(	499	));
			
 U508	: Somador_Exato_1 PORT MAP(
	A=> C(	572	),
	B=> E(	438	),
	Cin=> Carry( 	507	),
	Cout=> Carry( 	508	),
	S=> E(	500	));
			
 U509	: Somador_Exato_1 PORT MAP(
	A=> C(	573	),
	B=> E(	439	),
	Cin=> Carry( 	508	),
	Cout=> Carry( 	509	),
	S=> E(	501	));
			
 U510	: Somador_Exato_1 PORT MAP(
	A=> C(	574	),
	B=> E(	440	),
	Cin=> Carry( 	509	),
	Cout=> Carry( 	510	),
	S=> E(	502	));
			
 U511	: Somador_Exato_1 PORT MAP(
	A=> C(	575	),
	B=> Carry(	447	),
	Cin=> Carry( 	510	),
	Cout=> Carry( 	511	),
	S=> E(	503	));
---
			
 U512	: Somador_Exato_1 PORT MAP(
	A=> C(	576	),
	B=> E(	441	),
	Cin=> '0'	,
	Cout=> Carry( 	512	),
	S=> R(	9	));
			
 U513	: Somador_Exato_1 PORT MAP(
	A=> C(	577	),
	B=> E(	442	),
	Cin=> Carry( 	512	),
	Cout=> Carry( 	513	),
	S=> E(	504	));
			
 U514	: Somador_Exato_1 PORT MAP(
	A=> C(	578	),
	B=> E(	443	),
	Cin=> Carry( 	513	),
	Cout=> Carry( 	514	),
	S=> E(	505	));
			
 U515	: Somador_Exato_1 PORT MAP(
	A=> C(	579	),
	B=> E(	444	),
	Cin=> Carry( 	514	),
	Cout=> Carry( 	515	),
	S=> E(	506	));
			
 U516	: Somador_Exato_1 PORT MAP(
	A=> C(	580	),
	B=> E(	445	),
	Cin=> Carry( 	515	),
	Cout=> Carry( 	516	),
	S=> E(	507	));
			
 U517	: Somador_Exato_1 PORT MAP(
	A=> C(	581	),
	B=> E(	446	),
	Cin=> Carry( 	516	),
	Cout=> Carry( 	517	),
	S=> E(	508	));
			
 U518	: Somador_Exato_1 PORT MAP(
	A=> C(	582	),
	B=> E(	447	),
	Cin=> Carry( 	517	),
	Cout=> Carry( 	518	),
	S=> E(	509	));
			
 U519	: Somador_Exato_1 PORT MAP(
	A=> C(	583	),
	B=> E(	448	),
	Cin=> Carry( 	518	),
	Cout=> Carry( 	519	),
	S=> E(	510	));
			
 U520	: Somador_Exato_1 PORT MAP(
	A=> C(	584	),
	B=> E(	449	),
	Cin=> Carry( 	519	),
	Cout=> Carry( 	520	),
	S=> E(	511	));
			
 U521	: Somador_Exato_1 PORT MAP(
	A=> C(	585	),
	B=> E(	450	),
	Cin=> Carry( 	520	),
	Cout=> Carry( 	521	),
	S=> E(	512	));
			
 U522	: Somador_Exato_1 PORT MAP(
	A=> C(	586	),
	B=> E(	451	),
	Cin=> Carry( 	521	),
	Cout=> Carry( 	522	),
	S=> E(	513	));
			
 U523	: Somador_Exato_1 PORT MAP(
	A=> C(	587	),
	B=> E(	452	),
	Cin=> Carry( 	522	),
	Cout=> Carry( 	523	),
	S=> E(	514	));
			
 U524	: Somador_Exato_1 PORT MAP(
	A=> C(	588	),
	B=> E(	453	),
	Cin=> Carry( 	523	),
	Cout=> Carry( 	524	),
	S=> E(	515	));
			
 U525	: Somador_Exato_1 PORT MAP(
	A=> C(	589	),
	B=> E(	454	),
	Cin=> Carry( 	524	),
	Cout=> Carry( 	525	),
	S=> E(	516	));
			
 U526	: Somador_Exato_1 PORT MAP(
	A=> C(	590	),
	B=> E(	455	),
	Cin=> Carry( 	525	),
	Cout=> Carry( 	526	),
	S=> E(	517	));
			
 U527	: Somador_Exato_1 PORT MAP(
	A=> C(	591	),
	B=> E(	456	),
	Cin=> Carry( 	526	),
	Cout=> Carry( 	527	),
	S=> E(	518	));
			
 U528	: Somador_Exato_1 PORT MAP(
	A=> C(	592	),
	B=> E(	457	),
	Cin=> Carry( 	527	),
	Cout=> Carry( 	528	),
	S=> E(	519	));
			
 U529	: Somador_Exato_1 PORT MAP(
	A=> C(	593	),
	B=> E(	458	),
	Cin=> Carry( 	528	),
	Cout=> Carry( 	529	),
	S=> E(	520	));
			
 U530	: Somador_Exato_1 PORT MAP(
	A=> C(	594	),
	B=> E(	459	),
	Cin=> Carry( 	529	),
	Cout=> Carry( 	530	),
	S=> E(	521	));
			
 U531	: Somador_Exato_1 PORT MAP(
	A=> C(	595	),
	B=> E(	460	),
	Cin=> Carry( 	530	),
	Cout=> Carry( 	531	),
	S=> E(	522	));
			
 U532	: Somador_Exato_1 PORT MAP(
	A=> C(	596	),
	B=> E(	461	),
	Cin=> Carry( 	531	),
	Cout=> Carry( 	532	),
	S=> E(	523	));
			
 U533	: Somador_Exato_1 PORT MAP(
	A=> C(	597	),
	B=> E(	462	),
	Cin=> Carry( 	532	),
	Cout=> Carry( 	533	),
	S=> E(	524	));
			
 U534	: Somador_Exato_1 PORT MAP(
	A=> C(	598	),
	B=> E(	463	),
	Cin=> Carry( 	533	),
	Cout=> Carry( 	534	),
	S=> E(	525	));
			
 U535	: Somador_Exato_1 PORT MAP(
	A=> C(	599	),
	B=> E(	464	),
	Cin=> Carry( 	534	),
	Cout=> Carry( 	535	),
	S=> E(	526	));
			
 U536	: Somador_Exato_1 PORT MAP(
	A=> C(	600	),
	B=> E(	465	),
	Cin=> Carry( 	535	),
	Cout=> Carry( 	536	),
	S=> E(	527	));
			
 U537	: Somador_Exato_1 PORT MAP(
	A=> C(	601	),
	B=> E(	466	),
	Cin=> Carry( 	536	),
	Cout=> Carry( 	537	),
	S=> E(	528	));
			
 U538	: Somador_Exato_1 PORT MAP(
	A=> C(	602	),
	B=> E(	467	),
	Cin=> Carry( 	537	),
	Cout=> Carry( 	538	),
	S=> E(	529	));
			
 U539	: Somador_Exato_1 PORT MAP(
	A=> C(	603	),
	B=> E(	468	),
	Cin=> Carry( 	538	),
	Cout=> Carry( 	539	),
	S=> E(	530	));
			
 U540	: Somador_Exato_1 PORT MAP(
	A=> C(	604	),
	B=> E(	469	),
	Cin=> Carry( 	539	),
	Cout=> Carry( 	540	),
	S=> E(	531	));
			
 U541	: Somador_Exato_1 PORT MAP(
	A=> C(	605	),
	B=> E(	470	),
	Cin=> Carry( 	540	),
	Cout=> Carry( 	541	),
	S=> E(	532	));
			
 U542	: Somador_Exato_1 PORT MAP(
	A=> C(	606	),
	B=> E(	471	),
	Cin=> Carry( 	541	),
	Cout=> Carry( 	542	),
	S=> E(	533	));
			
 U543	: Somador_Exato_1 PORT MAP(
	A=> C(	607	),
	B=> E(	472	),
	Cin=> Carry( 	542	),
	Cout=> Carry( 	543	),
	S=> E(	534	));
			
 U544	: Somador_Exato_1 PORT MAP(
	A=> C(	608	),
	B=> E(	473	),
	Cin=> Carry( 	543	),
	Cout=> Carry( 	544	),
	S=> E(	535	));
			
 U545	: Somador_Exato_1 PORT MAP(
	A=> C(	609	),
	B=> E(	474	),
	Cin=> Carry( 	544	),
	Cout=> Carry( 	545	),
	S=> E(	536	));
			
 U546	: Somador_Exato_1 PORT MAP(
	A=> C(	610	),
	B=> E(	475	),
	Cin=> Carry( 	545	),
	Cout=> Carry( 	546	),
	S=> E(	537	));
			
 U547	: Somador_Exato_1 PORT MAP(
	A=> C(	611	),
	B=> E(	476	),
	Cin=> Carry( 	546	),
	Cout=> Carry( 	547	),
	S=> E(	538	));
			
 U548	: Somador_Exato_1 PORT MAP(
	A=> C(	612	),
	B=> E(	477	),
	Cin=> Carry( 	547	),
	Cout=> Carry( 	548	),
	S=> E(	539	));
 			
 U549	: Somador_Exato_1 PORT MAP(
	A=> C(	613	),
	B=> E(	478	),
	Cin=> Carry( 	548	),
	Cout=> Carry( 	549	),
	S=> E(	540	));
			
 U550	: Somador_Exato_1 PORT MAP(
	A=> C(	614	),
	B=> E(	479	),
	Cin=> Carry( 	549	),
	Cout=> Carry( 	550	),
	S=> E(	541	));
			
 U551	: Somador_Exato_1 PORT MAP(
	A=> C(	615	),
	B=> E(	480	),
	Cin=> Carry( 	550	),
	Cout=> Carry( 	551	),
	S=> E(	542	));
			
 U552	: Somador_Exato_1 PORT MAP(
	A=> C(	616	),
	B=> E(	481	),
	Cin=> Carry( 	551	),
	Cout=> Carry( 	552	),
	S=> E(	543	));
			
 U553	: Somador_Exato_1 PORT MAP(
	A=> C(	617	),
	B=> E(	482	),
	Cin=> Carry( 	552	),
	Cout=> Carry( 	553	),
	S=> E(	544	));
			
 U554	: Somador_Exato_1 PORT MAP(
	A=> C(	618	),
	B=> E(	483	),
	Cin=> Carry( 	553	),
	Cout=> Carry( 	554	),
	S=> E(	545	));
			
 U555	: Somador_Exato_1 PORT MAP(
	A=> C(	619	),
	B=> E(	484	),
	Cin=> Carry( 	554	),
	Cout=> Carry( 	555	),
	S=> E(	546	));
			
 U556	: Somador_Exato_1 PORT MAP(
	A=> C(	620	),
	B=> E(	485	),
	Cin=> Carry( 	555	),
	Cout=> Carry( 	556	),
	S=> E(	547	));
			
 U557	: Somador_Exato_1 PORT MAP(
	A=> C(	621	),
	B=> E(	486	),
	Cin=> Carry( 	556	),
	Cout=> Carry( 	557	),
	S=> E(	548	));
			
 U558	: Somador_Exato_1 PORT MAP(
	A=> C(	622	),
	B=> E(	487	),
	Cin=> Carry( 	557	),
	Cout=> Carry( 	558	),
	S=> E(	549	));
			
 U559	: Somador_Exato_1 PORT MAP(
	A=> C(	623	),
	B=> E(	488	),
	Cin=> Carry( 	558	),
	Cout=> Carry( 	559	),
	S=> E(	550	));
			
 U560	: Somador_Exato_1 PORT MAP(
	A=> C(	624	),
	B=> E(	489	),
	Cin=> Carry( 	559	),
	Cout=> Carry( 	560	),
	S=> E(	551	));
			
 U561	: Somador_Exato_1 PORT MAP(
	A=> C(	625	),
	B=> E(	490	),
	Cin=> Carry( 	560	),
	Cout=> Carry( 	561	),
	S=> E(	552	));
			
 U562	: Somador_Exato_1 PORT MAP(
	A=> C(	626	),
	B=> E(	491	),
	Cin=> Carry( 	561	),
	Cout=> Carry( 	562	),
	S=> E(	553	));
			
 U563	: Somador_Exato_1 PORT MAP(
	A=> C(	627	),
	B=> E(	492	),
	Cin=> Carry( 	562	),
	Cout=> Carry( 	563	),
	S=> E(	554	));
			
 U564	: Somador_Exato_1 PORT MAP(
	A=> C(	628	),
	B=> E(	493	),
	Cin=> Carry( 	563	),
	Cout=> Carry( 	564	),
	S=> E(	555	));
			
 U565	: Somador_Exato_1 PORT MAP(
	A=> C(	629	),
	B=> E(	494	),
	Cin=> Carry( 	564	),
	Cout=> Carry( 	565	),
	S=> E(	556	));
			
 U566	: Somador_Exato_1 PORT MAP(
	A=> C(	630	),
	B=> E(	495	),
	Cin=> Carry( 	565	),
	Cout=> Carry( 	566	),
	S=> E(	557	));
			
 U567	: Somador_Exato_1 PORT MAP(
	A=> C(	631	),
	B=> E(	496	),
	Cin=> Carry( 	566	),
	Cout=> Carry( 	567	),
	S=> E(	558	));
			
 U568	: Somador_Exato_1 PORT MAP(
	A=> C(	632	),
	B=> E(	497	),
	Cin=> Carry( 	567	),
	Cout=> Carry( 	568	),
	S=> E(	559	));
			
 U569	: Somador_Exato_1 PORT MAP(
	A=> C(	633	),
	B=> E(	498	),
	Cin=> Carry( 	568	),
	Cout=> Carry( 	569	),
	S=> E(	560	));
			
 U570	: Somador_Exato_1 PORT MAP(
	A=> C(	634	),
	B=> E(	499	),
	Cin=> Carry( 	569	),
	Cout=> Carry( 	570	),
	S=> E(	561	));
			
 U571	: Somador_Exato_1 PORT MAP(
	A=> C(	635	),
	B=> E(	500	),
	Cin=> Carry( 	570	),
	Cout=> Carry( 	571	),
	S=> E(	562	));
			
 U572	: Somador_Exato_1 PORT MAP(
	A=> C(	636	),
	B=> E(	501	),
	Cin=> Carry( 	571	),
	Cout=> Carry( 	572	),
	S=> E(	563	));
			
 U573	: Somador_Exato_1 PORT MAP(
	A=> C(	637	),
	B=> E(	502	),
	Cin=> Carry( 	572	),
	Cout=> Carry( 	573	),
	S=> E(	564	));
			
 U574	: Somador_Exato_1 PORT MAP(
	A=> C(	638	),
	B=> E(	503	),
	Cin=> Carry( 	573	),
	Cout=> Carry( 	574	),
	S=> E(	565	));
			
 U575	: Somador_Exato_1 PORT MAP(
	A => C(639),
	B => Carry(511),
	Cin => Carry(574),
	Cout => Carry(575),
	S => E(566));

			
 U576	: Somador_Exato_1 PORT MAP(
	A=> C(	640	),
	B=> E(	504	),
	Cin=> '0'	,
	Cout=> Carry( 	576	),
	S=> R(	10	));
			
 U577	: Somador_Exato_1 PORT MAP(
	A=> C(	641	),
	B=> E(	505	),
	Cin=> Carry( 	576	),
	Cout=> Carry( 	577	),
	S=> E(	567	));
			
 U578	: Somador_Exato_1 PORT MAP(
	A=> C(	642	),
	B=> E(	506	),
	Cin=> Carry( 	577	),
	Cout=> Carry( 	578	),
	S=> E(	568	));
			
 U579	: Somador_Exato_1 PORT MAP(
	A=> C(	643	),
	B=> E(	507	),
	Cin=> Carry( 	578	),
	Cout=> Carry( 	579	),
	S=> E(	569	));
			
 U580	: Somador_Exato_1 PORT MAP(
	A=> C(	644	),
	B=> E(	508	),
	Cin=> Carry( 	579	),
	Cout=> Carry( 	580	),
	S=> E(	570	));
			
 U581	: Somador_Exato_1 PORT MAP(
	A=> C(	645	),
	B=> E(	509	),
	Cin=> Carry( 	580	),
	Cout=> Carry( 	581	),
	S=> E(	571	));
			
 U582	: Somador_Exato_1 PORT MAP(
	A=> C(	646	),
	B=> E(	510	),
	Cin=> Carry( 	581	),
	Cout=> Carry( 	582	),
	S=> E(	572	));
			
 U583	: Somador_Exato_1 PORT MAP(
	A=> C(	647	),
	B=> E(	511	),
	Cin=> Carry( 	582	),
	Cout=> Carry( 	583	),
	S=> E(	573	));
			
 U584	: Somador_Exato_1 PORT MAP(
	A=> C(	648	),
	B=> E(	512	),
	Cin=> Carry( 	583	),
	Cout=> Carry( 	584	),
	S=> E(	574	));
			
 U585	: Somador_Exato_1 PORT MAP(
	A=> C(	649	),
	B=> E(	513	),
	Cin=> Carry( 	584	),
	Cout=> Carry( 	585	),
	S=> E(	575	));
			
 U586	: Somador_Exato_1 PORT MAP(
	A=> C(	650	),
	B=> E(	514	),
	Cin=> Carry( 	585	),
	Cout=> Carry( 	586	),
	S=> E(	576	));
			
 U587	: Somador_Exato_1 PORT MAP(
	A=> C(	651	),
	B=> E(	515	),
	Cin=> Carry( 	586	),
	Cout=> Carry( 	587	),
	S=> E(	577	));
			
 U588	: Somador_Exato_1 PORT MAP(
	A=> C(	652	),
	B=> E(	516	),
	Cin=> Carry( 	587	),
	Cout=> Carry( 	588	),
	S=> E(	578	));
			
 U589	: Somador_Exato_1 PORT MAP(
	A=> C(	653	),
	B=> E(	517	),
	Cin=> Carry( 	588	),
	Cout=> Carry( 	589	),
	S=> E(	579	));
			
 U590	: Somador_Exato_1 PORT MAP(
	A=> C(	654	),
	B=> E(	518	),
	Cin=> Carry( 	589	),
	Cout=> Carry( 	590	),
	S=> E(	580	));
			
 U591	: Somador_Exato_1 PORT MAP(
	A=> C(	655	),
	B=> E(	519	),
	Cin=> Carry( 	590	),
	Cout=> Carry( 	591	),
	S=> E(	581	));
			
 U592	: Somador_Exato_1 PORT MAP(
	A=> C(	656	),
	B=> E(	520	),
	Cin=> Carry( 	591	),
	Cout=> Carry( 	592	),
	S=> E(	582	));
			
 U593	: Somador_Exato_1 PORT MAP(
	A=> C(	657	),
	B=> E(	521	),
	Cin=> Carry( 	592	),
	Cout=> Carry( 	593	),
	S=> E(	583	));
			
 U594	: Somador_Exato_1 PORT MAP(
	A=> C(	658	),
	B=> E(	522	),
	Cin=> Carry( 	593	),
	Cout=> Carry( 	594	),
	S=> E(	584	));
			
 U595	: Somador_Exato_1 PORT MAP(
	A=> C(	659	),
	B=> E(	523	),
	Cin=> Carry( 	594	),
	Cout=> Carry( 	595	),
	S=> E(	585	));
			
 U596	: Somador_Exato_1 PORT MAP(
	A=> C(	660	),
	B=> E(	524	),
	Cin=> Carry( 	595	),
	Cout=> Carry( 	596	),
	S=> E(	586	));
			
 U597	: Somador_Exato_1 PORT MAP(
	A=> C(	661	),
	B=> E(	525	),
	Cin=> Carry( 	596	),
	Cout=> Carry( 	597	),
	S=> E(	587	));
			
 U598	: Somador_Exato_1 PORT MAP(
	A=> C(	662	),
	B=> E(	526	),
	Cin=> Carry( 	597	),
	Cout=> Carry( 	598	),
	S=> E(	588	));
			
 U599	: Somador_Exato_1 PORT MAP(
	A=> C(	663	),
	B=> E(	527	),
	Cin=> Carry( 	598	),
	Cout=> Carry( 	599	),
	S=> E(	589	));
			
 U600	: Somador_Exato_1 PORT MAP(
	A=> C(	664	),
	B=> E(	528	),
	Cin=> Carry( 	599	),
	Cout=> Carry( 	600	),
	S=> E(	590	));
			
 U601	: Somador_Exato_1 PORT MAP(
	A=> C(	665	),
	B=> E(	529	),
	Cin=> Carry( 	600	),
	Cout=> Carry( 	601	),
	S=> E(	591	));
			
 U602	: Somador_Exato_1 PORT MAP(
	A=> C(	666	),
	B=> E(	530	),
	Cin=> Carry( 	601	),
	Cout=> Carry( 	602	),
	S=> E(	592	));
			
 U603	: Somador_Exato_1 PORT MAP(
	A=> C(	667	),
	B=> E(	531	),
	Cin=> Carry( 	602	),
	Cout=> Carry( 	603	),
	S=> E(	593	));
			
 U604	: Somador_Exato_1 PORT MAP(
	A=> C(	668	),
	B=> E(	532	),
	Cin=> Carry( 	603	),
	Cout=> Carry( 	604	),
	S=> E(	594	));
			
 U605	: Somador_Exato_1 PORT MAP(
	A=> C(	669	),
	B=> E(	533	),
	Cin=> Carry( 	604	),
	Cout=> Carry( 	605	),
	S=> E(	595	));
			
 U606	: Somador_Exato_1 PORT MAP(
	A=> C(	670	),
	B=> E(	534	),
	Cin=> Carry( 	605	),
	Cout=> Carry( 	606	),
	S=> E(	596	));
			
 U607	: Somador_Exato_1 PORT MAP(
	A=> C(	671	),
	B=> E(	535	),
	Cin=> Carry( 	606	),
	Cout=> Carry( 	607	),
	S=> E(	597	));
			
 U608	: Somador_Exato_1 PORT MAP(
	A=> C(	672	),
	B=> E(	536	),
	Cin=> Carry( 	607	),
	Cout=> Carry( 	608	),
	S=> E(	598	));
			
 U609	: Somador_Exato_1 PORT MAP(
	A=> C(	673	),
	B=> E(	537	),
	Cin=> Carry( 	608	),
	Cout=> Carry( 	609	),
	S=> E(	599	));
			
 U610	: Somador_Exato_1 PORT MAP(
	A=> C(	674	),
	B=> E(	538	),
	Cin=> Carry( 	609	),
	Cout=> Carry( 	610	),
	S=> E(	600	));
			
 U611	: Somador_Exato_1 PORT MAP(
	A=> C(	675	),
	B=> E(	539	),
	Cin=> Carry( 	610	),
	Cout=> Carry( 	611	),
	S=> E(	601	));
			
 U612	: Somador_Exato_1 PORT MAP(
	A=> C(	676	),
	B=> E(	540	),
	Cin=> Carry( 	611	),
	Cout=> Carry( 	612	),
	S=> E(	602	));
			
 U613	: Somador_Exato_1 PORT MAP(
	A=> C(	677	),
	B=> E(	541	),
	Cin=> Carry( 	612	),
	Cout=> Carry( 	613	),
	S=> E(	603	));
			
 U614	: Somador_Exato_1 PORT MAP(
	A=> C(	678	),
	B=> E(	542	),
	Cin=> Carry( 	613	),
	Cout=> Carry( 	614	),
	S=> E(	604	));
			
 U615	: Somador_Exato_1 PORT MAP(
	A=> C(	679	),
	B=> E(	543	),
	Cin=> Carry( 	614	),
	Cout=> Carry( 	615	),
	S=> E(	605	));
			
 U616	: Somador_Exato_1 PORT MAP(
	A=> C(	680	),
	B=> E(	544	),
	Cin=> Carry( 	615	),
	Cout=> Carry( 	616	),
	S=> E(	606	));
			
 U617	: Somador_Exato_1 PORT MAP(
	A=> C(	681	),
	B=> E(	545	),
	Cin=> Carry( 	616	),
	Cout=> Carry( 	617	),
	S=> E(	607	));
			
 U618	: Somador_Exato_1 PORT MAP(
	A=> C(	682	),
	B=> E(	546	),
	Cin=> Carry( 	617	),
	Cout=> Carry( 	618	),
	S=> E(	608	));
			
 U619	: Somador_Exato_1 PORT MAP(
	A=> C(	683	),
	B=> E(	547	),
	Cin=> Carry( 	618	),
	Cout=> Carry( 	619	),
	S=> E(	609	));
			
 U620	: Somador_Exato_1 PORT MAP(
	A=> C(	684	),
	B=> E(	548	),
	Cin=> Carry( 	619	),
	Cout=> Carry( 	620	),
	S=> E(	610	));
			
 U621	: Somador_Exato_1 PORT MAP(
	A=> C(	685	),
	B=> E(	549	),
	Cin=> Carry( 	620	),
	Cout=> Carry( 	621	),
	S=> E(	611	));
			
 U622	: Somador_Exato_1 PORT MAP(
	A=> C(	686	),
	B=> E(	550	),
	Cin=> Carry( 	621	),
	Cout=> Carry( 	622	),
	S=> E(	612	));
			
 U623	: Somador_Exato_1 PORT MAP(
	A=> C(	687	),
	B=> E(	551	),
	Cin=> Carry( 	622	),
	Cout=> Carry( 	623	),
	S=> E(	613	));
			
 U624	: Somador_Exato_1 PORT MAP(
	A=> C(	688	),
	B=> E(	552	),
	Cin=> Carry( 	623	),
	Cout=> Carry( 	624	),
	S=> E(	614	));
			
 U625	: Somador_Exato_1 PORT MAP(
	A=> C(	689	),
	B=> E(	553	),
	Cin=> Carry( 	624	),
	Cout=> Carry( 	625	),
	S=> E(	615	));
			
 U626	: Somador_Exato_1 PORT MAP(
	A=> C(	690	),
	B=> E(	554	),
	Cin=> Carry( 	625	),
	Cout=> Carry( 	626	),
	S=> E(	616	));
			
 U627	: Somador_Exato_1 PORT MAP(
	A=> C(	691	),
	B=> E(	555	),
	Cin=> Carry( 	626	),
	Cout=> Carry( 	627	),
	S=> E(	617	));
			
 U628	: Somador_Exato_1 PORT MAP(
	A=> C(	692	),
	B=> E(	556	),
	Cin=> Carry( 	627	),
	Cout=> Carry( 	628	),
	S=> E(	618	));
			
 U629	: Somador_Exato_1 PORT MAP(
	A=> C(	693	),
	B=> E(	557	),
	Cin=> Carry( 	628	),
	Cout=> Carry( 	629	),
	S=> E(	619	));
			
 U630	: Somador_Exato_1 PORT MAP(
	A=> C(	694	),
	B=> E(	558	),
	Cin=> Carry( 	629	),
	Cout=> Carry( 	630	),
	S=> E(	620	));
			
 U631	: Somador_Exato_1 PORT MAP(
	A=> C(	695	),
	B=> E(	559	),
	Cin=> Carry( 	630	),
	Cout=> Carry( 	631	),
	S=> E(	621	));
			
 U632	: Somador_Exato_1 PORT MAP(
	A=> C(	696	),
	B=> E(	560	),
	Cin=> Carry( 	631	),
	Cout=> Carry( 	632	),
	S=> E(	622	));
			
 U633	: Somador_Exato_1 PORT MAP(
	A=> C(	697	),
	B=> E(	561	),
	Cin=> Carry( 	632	),
	Cout=> Carry( 	633	),
	S=> E(	623	));
			
 U634	: Somador_Exato_1 PORT MAP(
	A=> C(	698	),
	B=> E(	562	),
	Cin=> Carry( 	633	),
	Cout=> Carry( 	634	),
	S=> E(	624	));
			
 U635	: Somador_Exato_1 PORT MAP(
	A=> C(	699	),
	B=> E(	563	),
	Cin=> Carry( 	634	),
	Cout=> Carry( 	635	),
	S=> E(	625	));
			
 U636	: Somador_Exato_1 PORT MAP(
	A=> C(	700	),
	B=> E(	564	),
	Cin=> Carry( 	635	),
	Cout=> Carry( 	636	),
	S=> E(	626	));
			
 U637	: Somador_Exato_1 PORT MAP(
	A=> C(	701	),
	B=> E(	565	),
	Cin=> Carry( 	636	),
	Cout=> Carry( 	637	),
	S=> E(	627	));
			
 U638	: Somador_Exato_1 PORT MAP(
	A=> C(	702	),
	B=> E(	566	),
	Cin=> Carry( 	637	),
	Cout=> Carry( 	638	),
	S=> E(	628	));
			
 U639	: Somador_Exato_1 PORT MAP(
	A=> C(	703	),
	B=> Carry(	575	),
	Cin=> Carry( 	638	),
	Cout=> Carry( 	639	),
	S=> E(	629	));

			
 U640	: Somador_Exato_1 PORT MAP(
	A=> C(	704	),
	B=> E(	567	),
	Cin=> '0'	,
	Cout=> Carry( 	640	),
	S=> R(	11	));
			
 U641	: Somador_Exato_1 PORT MAP(
	A=> C(	705	),
	B=> E(	568	),
	Cin=> Carry( 	640	),
	Cout=> Carry( 	641	),
	S=> E(	630	));
			
 U642	: Somador_Exato_1 PORT MAP(
	A=> C(	706	),
	B=> E(	569	),
	Cin=> Carry( 	641	),
	Cout=> Carry( 	642	),
	S=> E(	631	));
			
 U643	: Somador_Exato_1 PORT MAP(
	A=> C(	707	),
	B=> E(	570	),
	Cin=> Carry( 	642	),
	Cout=> Carry( 	643	),
	S=> E(	632	));
			
 U644	: Somador_Exato_1 PORT MAP(
	A=> C(	708	),
	B=> E(	571	),
	Cin=> Carry( 	643	),
	Cout=> Carry( 	644	),
	S=> E(	633	));
			
 U645	: Somador_Exato_1 PORT MAP(
	A=> C(	709	),
	B=> E(	572	),
	Cin=> Carry( 	644	),
	Cout=> Carry( 	645	),
	S=> E(	634	));
			
 U646	: Somador_Exato_1 PORT MAP(
	A=> C(	710	),
	B=> E(	573	),
	Cin=> Carry( 	645	),
	Cout=> Carry( 	646	),
	S=> E(	635	));
			
 U647	: Somador_Exato_1 PORT MAP(
	A=> C(	711	),
	B=> E(	574	),
	Cin=> Carry( 	646	),
	Cout=> Carry( 	647	),
	S=> E(	636	));
			
 U648	: Somador_Exato_1 PORT MAP(
	A=> C(	712	),
	B=> E(	575	),
	Cin=> Carry( 	647	),
	Cout=> Carry( 	648	),
	S=> E(	637	));
			
 U649	: Somador_Exato_1 PORT MAP(
	A=> C(	713	),
	B=> E(	576	),
	Cin=> Carry( 	648	),
	Cout=> Carry( 	649	),
	S=> E(	638	));
			
 U650	: Somador_Exato_1 PORT MAP(
	A=> C(	714	),
	B=> E(	577	),
	Cin=> Carry( 	649	),
	Cout=> Carry( 	650	),
	S=> E(	639	));
			
 U651	: Somador_Exato_1 PORT MAP(
	A=> C(	715	),
	B=> E(	578	),
	Cin=> Carry( 	650	),
	Cout=> Carry( 	651	),
	S=> E(	640	));
			
 U652	: Somador_Exato_1 PORT MAP(
	A=> C(	716	),
	B=> E(	579	),
	Cin=> Carry( 	651	),
	Cout=> Carry( 	652	),
	S=> E(	641	));
			
 U653	: Somador_Exato_1 PORT MAP(
	A=> C(	717	),
	B=> E(	580	),
	Cin=> Carry( 	652	),
	Cout=> Carry( 	653	),
	S=> E(	642	));
			
 U654	: Somador_Exato_1 PORT MAP(
	A=> C(	718	),
	B=> E(	581	),
	Cin=> Carry( 	653	),
	Cout=> Carry( 	654	),
	S=> E(	643	));
			
 U655	: Somador_Exato_1 PORT MAP(
	A=> C(	719	),
	B=> E(	582	),
	Cin=> Carry( 	654	),
	Cout=> Carry( 	655	),
	S=> E(	644	));
			
 U656	: Somador_Exato_1 PORT MAP(
	A=> C(	720	),
	B=> E(	583	),
	Cin=> Carry( 	655	),
	Cout=> Carry( 	656	),
	S=> E(	645	));
			
 U657	: Somador_Exato_1 PORT MAP(
	A=> C(	721	),
	B=> E(	584	),
	Cin=> Carry( 	656	),
	Cout=> Carry( 	657	),
	S=> E(	646	));
			
 U658	: Somador_Exato_1 PORT MAP(
	A=> C(	722	),
	B=> E(	585	),
	Cin=> Carry( 	657	),
	Cout=> Carry( 	658	),
	S=> E(	647	));
			
 U659	: Somador_Exato_1 PORT MAP(
	A=> C(	723	),
	B=> E(	586	),
	Cin=> Carry( 	658	),
	Cout=> Carry( 	659	),
	S=> E(	648	));
			
 U660	: Somador_Exato_1 PORT MAP(
	A=> C(	724	),
	B=> E(	587	),
	Cin=> Carry( 	659	),
	Cout=> Carry( 	660	),
	S=> E(	649	));
			
 U661	: Somador_Exato_1 PORT MAP(
	A=> C(	725	),
	B=> E(	588	),
	Cin=> Carry( 	660	),
	Cout=> Carry( 	661	),
	S=> E(	650	));
			
 U662	: Somador_Exato_1 PORT MAP(
	A=> C(	726	),
	B=> E(	589	),
	Cin=> Carry( 	661	),
	Cout=> Carry( 	662	),
	S=> E(	651	));
			
 U663	: Somador_Exato_1 PORT MAP(
	A=> C(	727	),
	B=> E(	590	),
	Cin=> Carry( 	662	),
	Cout=> Carry( 	663	),
	S=> E(	652	));
			
 U664	: Somador_Exato_1 PORT MAP(
	A=> C(	728	),
	B=> E(	591	),
	Cin=> Carry( 	663	),
	Cout=> Carry( 	664	),
	S=> E(	653	));
			
 U665	: Somador_Exato_1 PORT MAP(
	A=> C(	729	),
	B=> E(	592	),
	Cin=> Carry( 	664	),
	Cout=> Carry( 	665	),
	S=> E(	654	));
			
 U666	: Somador_Exato_1 PORT MAP(
	A=> C(	730	),
	B=> E(	593	),
	Cin=> Carry( 	665	),
	Cout=> Carry( 	666	),
	S=> E(	655	));
			
 U667	: Somador_Exato_1 PORT MAP(
	A=> C(	731	),
	B=> E(	594	),
	Cin=> Carry( 	666	),
	Cout=> Carry( 	667	),
	S=> E(	656	));
			
 U668	: Somador_Exato_1 PORT MAP(
	A=> C(	732	),
	B=> E(	595	),
	Cin=> Carry( 	667	),
	Cout=> Carry( 	668	),
	S=> E(	657	));
			
 U669	: Somador_Exato_1 PORT MAP(
	A=> C(	733	),
	B=> E(	596	),
	Cin=> Carry( 	668	),
	Cout=> Carry( 	669	),
	S=> E(	658	));
			
 U670	: Somador_Exato_1 PORT MAP(
	A=> C(	734	),
	B=> E(	597	),
	Cin=> Carry( 	669	),
	Cout=> Carry( 	670	),
	S=> E(	659	));
			
 U671	: Somador_Exato_1 PORT MAP(
	A=> C(	735	),
	B=> E(	598	),
	Cin=> Carry( 	670	),
	Cout=> Carry( 	671	),
	S=> E(	660	));
			
 U672	: Somador_Exato_1 PORT MAP(
	A=> C(	736	),
	B=> E(	599	),
	Cin=> Carry( 	671	),
	Cout=> Carry( 	672	),
	S=> E(	661	));
			
 U673	: Somador_Exato_1 PORT MAP(
	A=> C(	737	),
	B=> E(	600	),
	Cin=> Carry( 	672	),
	Cout=> Carry( 	673	),
	S=> E(	662	));
			
 U674	: Somador_Exato_1 PORT MAP(
	A=> C(	738	),
	B=> E(	601	),
	Cin=> Carry( 	673	),
	Cout=> Carry( 	674	),
	S=> E(	663	));
			
 U675	: Somador_Exato_1 PORT MAP(
	A=> C(	739	),
	B=> E(	602	),
	Cin=> Carry( 	674	),
	Cout=> Carry( 	675	),
	S=> E(	664	));
			
 U676	: Somador_Exato_1 PORT MAP(
	A=> C(	740	),
	B=> E(	603	),
	Cin=> Carry( 	675	),
	Cout=> Carry( 	676	),
	S=> E(	665	));
			
 U677	: Somador_Exato_1 PORT MAP(
	A=> C(	741	),
	B=> E(	604	),
	Cin=> Carry( 	676	),
	Cout=> Carry( 	677	),
	S=> E(	666	));
			
 U678	: Somador_Exato_1 PORT MAP(
	A=> C(	742	),
	B=> E(	605	),
	Cin=> Carry( 	677	),
	Cout=> Carry( 	678	),
	S=> E(	667	));
			
 U679	: Somador_Exato_1 PORT MAP(
	A=> C(	743	),
	B=> E(	606	),
	Cin=> Carry( 	678	),
	Cout=> Carry( 	679	),
	S=> E(	668	));
			
 U680	: Somador_Exato_1 PORT MAP(
	A=> C(	744	),
	B=> E(	607	),
	Cin=> Carry( 	679	),
	Cout=> Carry( 	680	),
	S=> E(	669	));
			
 U681	: Somador_Exato_1 PORT MAP(
	A=> C(	745	),
	B=> E(	608	),
	Cin=> Carry( 	680	),
	Cout=> Carry( 	681	),
	S=> E(	670	));
			
 U682	: Somador_Exato_1 PORT MAP(
	A=> C(	746	),
	B=> E(	609	),
	Cin=> Carry( 	681	),
	Cout=> Carry( 	682	),
	S=> E(	671	));
			
 U683	: Somador_Exato_1 PORT MAP(
	A=> C(	747	),
	B=> E(	610	),
	Cin=> Carry( 	682	),
	Cout=> Carry( 	683	),
	S=> E(	672	));
			
 U684	: Somador_Exato_1 PORT MAP(
	A=> C(	748	),
	B=> E(	611	),
	Cin=> Carry( 	683	),
	Cout=> Carry( 	684	),
	S=> E(	673	));
			
 U685	: Somador_Exato_1 PORT MAP(
	A=> C(	749	),
	B=> E(	612	),
	Cin=> Carry( 	684	),
	Cout=> Carry( 	685	),
	S=> E(	674	));
			
 U686	: Somador_Exato_1 PORT MAP(
	A=> C(	750	),
	B=> E(	613	),
	Cin=> Carry( 	685	),
	Cout=> Carry( 	686	),
	S=> E(	675	));
			
 U687	: Somador_Exato_1 PORT MAP(
	A=> C(	751	),
	B=> E(	614	),
	Cin=> Carry( 	686	),
	Cout=> Carry( 	687	),
	S=> E(	676	));
			
 U688	: Somador_Exato_1 PORT MAP(
	A=> C(	752	),
	B=> E(	615	),
	Cin=> Carry( 	687	),
	Cout=> Carry( 	688	),
	S=> E(	677	));
			
 U689	: Somador_Exato_1 PORT MAP(
	A=> C(	753	),
	B=> E(	616	),
	Cin=> Carry( 	688	),
	Cout=> Carry( 	689	),
	S=> E(	678	));
			
 U690	: Somador_Exato_1 PORT MAP(
	A=> C(	754	),
	B=> E(	617	),
	Cin=> Carry( 	689	),
	Cout=> Carry( 	690	),
	S=> E(	679	));
			
 U691	: Somador_Exato_1 PORT MAP(
	A=> C(	755	),
	B=> E(	618	),
	Cin=> Carry( 	690	),
	Cout=> Carry( 	691	),
	S=> E(	680	));
			
 U692	: Somador_Exato_1 PORT MAP(
	A=> C(	756	),
	B=> E(	619	),
	Cin=> Carry( 	691	),
	Cout=> Carry( 	692	),
	S=> E(	681	));
			
 U693	: Somador_Exato_1 PORT MAP(
	A=> C(	757	),
	B=> E(	620	),
	Cin=> Carry( 	692	),
	Cout=> Carry( 	693	),
	S=> E(	682	));
			
 U694	: Somador_Exato_1 PORT MAP(
	A=> C(	758	),
	B=> E(	621	),
	Cin=> Carry( 	693	),
	Cout=> Carry( 	694	),
	S=> E(	683	));
			
 U695	: Somador_Exato_1 PORT MAP(
	A=> C(	759	),
	B=> E(	622	),
	Cin=> Carry( 	694	),
	Cout=> Carry( 	695	),
	S=> E(	684	));
			
 U696	: Somador_Exato_1 PORT MAP(
	A=> C(	760	),
	B=> E(	623	),
	Cin=> Carry( 	695	),
	Cout=> Carry( 	696	),
	S=> E(	685	));
			
 U697	: Somador_Exato_1 PORT MAP(
	A=> C(	761	),
	B=> E(	624	),
	Cin=> Carry( 	696	),
	Cout=> Carry( 	697	),
	S=> E(	686	));
			
 U698	: Somador_Exato_1 PORT MAP(
	A=> C(	762	),
	B=> E(	625	),
	Cin=> Carry( 	697	),
	Cout=> Carry( 	698	),
	S=> E(	687	));
			
 U699	: Somador_Exato_1 PORT MAP(
	A=> C(	763	),
	B=> E(	626	),
	Cin=> Carry( 	698	),
	Cout=> Carry( 	699	),
	S=> E(	688	));
			
 U700	: Somador_Exato_1 PORT MAP(
	A=> C(	764	),
	B=> E(	627	),
	Cin=> Carry( 	699	),
	Cout=> Carry( 	700	),
	S=> E(	689	));
			
 U701	: Somador_Exato_1 PORT MAP(
	A=> C(	765	),
	B=> E(	628	),
	Cin=> Carry( 	700	),
	Cout=> Carry( 	701	),
	S=> E(	690	));
			
 U702	: Somador_Exato_1 PORT MAP(
	A=> C(	766	),
	B=> E(	629	),
	Cin=> Carry( 	701	),
	Cout=> Carry( 	702	),
	S=> E(	691	));
			
 U703	: Somador_Exato_1 PORT MAP(
	A=> C(	767	),
	B=> Carry(	639	),
	Cin=> Carry( 	702	),
	Cout=> Carry( 	703	),
	S=> E(	692	));

			
 U704	: Somador_Exato_1 PORT MAP(
	A=> C(	768	),
	B=> E(	630	),
	Cin=> '0',
	Cout=> Carry( 	704	),
	S=> R(	12	));
			
 U705	: Somador_Exato_1 PORT MAP(
	A=> C(	769	),
	B=> E(	631	),
	Cin=> Carry( 	704	),
	Cout=> Carry( 	705	),
	S=> E(	693	));
			
 U706	: Somador_Exato_1 PORT MAP(
	A=> C(	770	),
	B=> E(	632	),
	Cin=> Carry( 	705	),
	Cout=> Carry( 	706	),
	S=> E(	694	));
			
 U707	: Somador_Exato_1 PORT MAP(
	A=> C(	771	),
	B=> E(	633	),
	Cin=> Carry( 	706	),
	Cout=> Carry( 	707	),
	S=> E(	695	));
			
 U708	: Somador_Exato_1 PORT MAP(
	A=> C(	772	),
	B=> E(	634	),
	Cin=> Carry( 	707	),
	Cout=> Carry( 	708	),
	S=> E(	696	));
			
 U709	: Somador_Exato_1 PORT MAP(
	A=> C(	773	),
	B=> E(	635	),
	Cin=> Carry( 	708	),
	Cout=> Carry( 	709	),
	S=> E(	697	));
			
 U710	: Somador_Exato_1 PORT MAP(
	A=> C(	774	),
	B=> E(	636	),
	Cin=> Carry( 	709	),
	Cout=> Carry( 	710	),
	S=> E(	698	));
			
 U711	: Somador_Exato_1 PORT MAP(
	A=> C(	775	),
	B=> E(	637	),
	Cin=> Carry( 	710	),
	Cout=> Carry( 	711	),
	S=> E(	699	));
			
 U712	: Somador_Exato_1 PORT MAP(
	A=> C(	776	),
	B=> E(	638	),
	Cin=> Carry( 	711	),
	Cout=> Carry( 	712	),
	S=> E(	700	));
			
 U713	: Somador_Exato_1 PORT MAP(
	A=> C(	777	),
	B=> E(	639	),
	Cin=> Carry( 	712	),
	Cout=> Carry( 	713	),
	S=> E(	701	));
			
 U714	: Somador_Exato_1 PORT MAP(
	A=> C(	778	),
	B=> E(	640	),
	Cin=> Carry( 	713	),
	Cout=> Carry( 	714	),
	S=> E(	702	));
			
 U715	: Somador_Exato_1 PORT MAP(
	A=> C(	779	),
	B=> E(	641	),
	Cin=> Carry( 	714	),
	Cout=> Carry( 	715	),
	S=> E(	703	));
			
 U716	: Somador_Exato_1 PORT MAP(
	A=> C(	780	),
	B=> E(	642	),
	Cin=> Carry( 	715	),
	Cout=> Carry( 	716	),
	S=> E(	704	));
			
 U717	: Somador_Exato_1 PORT MAP(
	A=> C(	781	),
	B=> E(	643	),
	Cin=> Carry( 	716	),
	Cout=> Carry( 	717	),
	S=> E(	705	));
			
 U718	: Somador_Exato_1 PORT MAP(
	A=> C(	782	),
	B=> E(	644	),
	Cin=> Carry( 	717	),
	Cout=> Carry( 	718	),
	S=> E(	706	));
			
 U719	: Somador_Exato_1 PORT MAP(
	A=> C(	783	),
	B=> E(	645	),
	Cin=> Carry( 	718	),
	Cout=> Carry( 	719	),
	S=> E(	707	));
			
 U720	: Somador_Exato_1 PORT MAP(
	A=> C(	784	),
	B=> E(	646	),
	Cin=> Carry( 	719	),
	Cout=> Carry( 	720	),
	S=> E(	708	));
			
 U721	: Somador_Exato_1 PORT MAP(
	A=> C(	785	),
	B=> E(	647	),
	Cin=> Carry( 	720	),
	Cout=> Carry( 	721	),
	S=> E(	709	));
			
 U722	: Somador_Exato_1 PORT MAP(
	A=> C(	786	),
	B=> E(	648	),
	Cin=> Carry( 	721	),
	Cout=> Carry( 	722	),
	S=> E(	710	));
			
 U723	: Somador_Exato_1 PORT MAP(
	A=> C(	787	),
	B=> E(	649	),
	Cin=> Carry( 	722	),
	Cout=> Carry( 	723	),
	S=> E(	711	));
			
 U724	: Somador_Exato_1 PORT MAP(
	A=> C(	788	),
	B=> E(	650	),
	Cin=> Carry( 	723	),
	Cout=> Carry( 	724	),
	S=> E(	712	));
			
 U725	: Somador_Exato_1 PORT MAP(
	A=> C(	789	),
	B=> E(	651	),
	Cin=> Carry( 	724	),
	Cout=> Carry( 	725	),
	S=> E(	713	));
			
 U726	: Somador_Exato_1 PORT MAP(
	A=> C(	790	),
	B=> E(	652	),
	Cin=> Carry( 	725	),
	Cout=> Carry( 	726	),
	S=> E(	714	));
			
 U727	: Somador_Exato_1 PORT MAP(
	A=> C(	791	),
	B=> E(	653	),
	Cin=> Carry( 	726	),
	Cout=> Carry( 	727	),
	S=> E(	715	));
			
 U728	: Somador_Exato_1 PORT MAP(
	A=> C(	792	),
	B=> E(	654	),
	Cin=> Carry( 	727	),
	Cout=> Carry( 	728	),
	S=> E(	716	));
			
 U729	: Somador_Exato_1 PORT MAP(
	A=> C(	793	),
	B=> E(	655	),
	Cin=> Carry( 	728	),
	Cout=> Carry( 	729	),
	S=> E(	717	));
			
 U730	: Somador_Exato_1 PORT MAP(
	A=> C(	794	),
	B=> E(	656	),
	Cin=> Carry( 	729	),
	Cout=> Carry( 	730	),
	S=> E(	718	));
			
 U731	: Somador_Exato_1 PORT MAP(
	A=> C(	795	),
	B=> E(	657	),
	Cin=> Carry( 	730	),
	Cout=> Carry( 	731	),
	S=> E(	719	));
			
 U732	: Somador_Exato_1 PORT MAP(
	A=> C(	796	),
	B=> E(	658	),
	Cin=> Carry( 	731	),
	Cout=> Carry( 	732	),
	S=> E(	720	));
			
 U733	: Somador_Exato_1 PORT MAP(
	A=> C(	797	),
	B=> E(	659	),
	Cin=> Carry( 	732	),
	Cout=> Carry( 	733	),
	S=> E(	721	));
			
 U734	: Somador_Exato_1 PORT MAP(
	A=> C(	798	),
	B=> E(	660	),
	Cin=> Carry( 	733	),
	Cout=> Carry( 	734	),
	S=> E(	722	));
			
 U735	: Somador_Exato_1 PORT MAP(
	A=> C(	799	),
	B=> E(	661	),
	Cin=> Carry( 	734	),
	Cout=> Carry( 	735	),
	S=> E(	723	));
			
 U736	: Somador_Exato_1 PORT MAP(
	A=> C(	800	),
	B=> E(	662	),
	Cin=> Carry( 	735	),
	Cout=> Carry( 	736	),
	S=> E(	724	));
			
 U737	: Somador_Exato_1 PORT MAP(
	A=> C(	801	),
	B=> E(	663	),
	Cin=> Carry( 	736	),
	Cout=> Carry( 	737	),
	S=> E(	725	));
			
 U738	: Somador_Exato_1 PORT MAP(
	A=> C(	802	),
	B=> E(	664	),
	Cin=> Carry( 	737	),
	Cout=> Carry( 	738	),
	S=> E(	726	));
			
 U739	: Somador_Exato_1 PORT MAP(
	A=> C(	803	),
	B=> E(	665	),
	Cin=> Carry( 	738	),
	Cout=> Carry( 	739	),
	S=> E(	727	));
			
 U740	: Somador_Exato_1 PORT MAP(
	A=> C(	804	),
	B=> E(	666	),
	Cin=> Carry( 	739	),
	Cout=> Carry( 	740	),
	S=> E(	728	));
			
 U741	: Somador_Exato_1 PORT MAP(
	A=> C(	805	),
	B=> E(	667	),
	Cin=> Carry( 	740	),
	Cout=> Carry( 	741	),
	S=> E(	729	));
			
 U742	: Somador_Exato_1 PORT MAP(
	A=> C(	806	),
	B=> E(	668	),
	Cin=> Carry( 	741	),
	Cout=> Carry( 	742	),
	S=> E(	730	));
			
 U743	: Somador_Exato_1 PORT MAP(
	A=> C(	807	),
	B=> E(	669	),
	Cin=> Carry( 	742	),
	Cout=> Carry( 	743	),
	S=> E(	731	));
			
 U744	: Somador_Exato_1 PORT MAP(
	A=> C(	808	),
	B=> E(	670	),
	Cin=> Carry( 	743	),
	Cout=> Carry( 	744	),
	S=> E(	732	));
			
 U745	: Somador_Exato_1 PORT MAP(
	A=> C(	809	),
	B=> E(	671	),
	Cin=> Carry( 	744	),
	Cout=> Carry( 	745	),
	S=> E(	733	));
			
 U746	: Somador_Exato_1 PORT MAP(
	A=> C(	810	),
	B=> E(	672	),
	Cin=> Carry( 	745	),
	Cout=> Carry( 	746	),
	S=> E(	734	));
			
 U747	: Somador_Exato_1 PORT MAP(
	A=> C(	811	),
	B=> E(	673	),
	Cin=> Carry( 	746	),
	Cout=> Carry( 	747	),
	S=> E(	735	));
			
 U748	: Somador_Exato_1 PORT MAP(
	A=> C(	812	),
	B=> E(	674	),
	Cin=> Carry( 	747	),
	Cout=> Carry( 	748	),
	S=> E(	736	));
			
 U749	: Somador_Exato_1 PORT MAP(
	A=> C(	813	),
	B=> E(	675	),
	Cin=> Carry( 	748	),
	Cout=> Carry( 	749	),
	S=> E(	737	));
			
 U750	: Somador_Exato_1 PORT MAP(
	A=> C(	814	),
	B=> E(	676	),
	Cin=> Carry( 	749	),
	Cout=> Carry( 	750	),
	S=> E(	738	));
			
 U751	: Somador_Exato_1 PORT MAP(
	A=> C(	815	),
	B=> E(	677	),
	Cin=> Carry( 	750	),
	Cout=> Carry( 	751	),
	S=> E(	739	));
			
 U752	: Somador_Exato_1 PORT MAP(
	A=> C(	816	),
	B=> E(	678	),
	Cin=> Carry( 	751	),
	Cout=> Carry( 	752	),
	S=> E(	740	));
			
 U753	: Somador_Exato_1 PORT MAP(
	A=> C(	817	),
	B=> E(	679	),
	Cin=> Carry( 	752	),
	Cout=> Carry( 	753	),
	S=> E(	741	));
			
 U754	: Somador_Exato_1 PORT MAP(
	A=> C(	818	),
	B=> E(	680	),
	Cin=> Carry( 	753	),
	Cout=> Carry( 	754	),
	S=> E(	742	));
			
 U755	: Somador_Exato_1 PORT MAP(
	A=> C(	819	),
	B=> E(	681	),
	Cin=> Carry( 	754	),
	Cout=> Carry( 	755	),
	S=> E(	743	));
			
 U756	: Somador_Exato_1 PORT MAP(
	A=> C(	820	),
	B=> E(	682	),
	Cin=> Carry( 	755	),
	Cout=> Carry( 	756	),
	S=> E(	744	));
			
 U757	: Somador_Exato_1 PORT MAP(
	A=> C(	821	),
	B=> E(	683	),
	Cin=> Carry( 	756	),
	Cout=> Carry( 	757	),
	S=> E(	745	));
			
 U758	: Somador_Exato_1 PORT MAP(
	A=> C(	822	),
	B=> E(	684	),
	Cin=> Carry( 	757	),
	Cout=> Carry( 	758	),
	S=> E(	746	));
			
 U759	: Somador_Exato_1 PORT MAP(
	A=> C(	823	),
	B=> E(	685	),
	Cin=> Carry( 	758	),
	Cout=> Carry( 	759	),
	S=> E(	747	));
			
 U760	: Somador_Exato_1 PORT MAP(
	A=> C(	824	),
	B=> E(	686	),
	Cin=> Carry( 	759	),
	Cout=> Carry( 	760	),
	S=> E(	748	));
			
 U761	: Somador_Exato_1 PORT MAP(
	A=> C(	825	),
	B=> E(	687	),
	Cin=> Carry( 	760	),
	Cout=> Carry( 	761	),
	S=> E(	749	));
			
 U762	: Somador_Exato_1 PORT MAP(
	A=> C(	826	),
	B=> E(	688	),
	Cin=> Carry( 	761	),
	Cout=> Carry( 	762	),
	S=> E(	750	));
			
 U763	: Somador_Exato_1 PORT MAP(
	A=> C(	827	),
	B=> E(	689	),
	Cin=> Carry( 	762	),
	Cout=> Carry( 	763	),
	S=> E(	751	));
			
 U764	: Somador_Exato_1 PORT MAP(
	A=> C(	828	),
	B=> E(	690	),
	Cin=> Carry( 	763	),
	Cout=> Carry( 	764	),
	S=> E(	752	));
			
 U765	: Somador_Exato_1 PORT MAP(
	A=> C(	829	),
	B=> E(	691	),
	Cin=> Carry( 	764	),
	Cout=> Carry( 	765	),
	S=> E(	753	));
			
 U766	: Somador_Exato_1 PORT MAP(
	A=> C(	830	),
	B=> E(	692	),
	Cin=> Carry( 	765	),
	Cout=> Carry( 	766	),
	S=> E(	754	));
			
 U767	: Somador_Exato_1 PORT MAP(
	A=> C(	831	),
	B=> Carry(	703	),
	Cin=> Carry( 	766	),
	Cout=> Carry( 	767	),
	S=> E(	755	));

			
 U768	: Somador_Exato_1 PORT MAP(
	A=> C(	832	),
	B=> E(	693	),
	Cin=> '0'	,
	Cout=> Carry( 	768	),
	S=> R(	13	));
			
 U769	: Somador_Exato_1 PORT MAP(
	A=> C(	833	),
	B=> E(	694	),
	Cin=> Carry( 	768	),
	Cout=> Carry( 	769	),
	S=> E(	756	));
			
 U770	: Somador_Exato_1 PORT MAP(
	A=> C(	834	),
	B=> E(	695	),
	Cin=> Carry( 	769	),
	Cout=> Carry( 	770	),
	S=> E(	757	));
			
 U771	: Somador_Exato_1 PORT MAP(
	A=> C(	835	),
	B=> E(	696	),
	Cin=> Carry( 	770	),
	Cout=> Carry( 	771	),
	S=> E(	758	));
			
 U772	: Somador_Exato_1 PORT MAP(
	A=> C(	836	),
	B=> E(	697	),
	Cin=> Carry( 	771	),
	Cout=> Carry( 	772	),
	S=> E(	759	));
			
 U773	: Somador_Exato_1 PORT MAP(
	A=> C(	837	),
	B=> E(	698	),
	Cin=> Carry( 	772	),
	Cout=> Carry( 	773	),
	S=> E(	760	));
			
 U774	: Somador_Exato_1 PORT MAP(
	A=> C(	838	),
	B=> E(	699	),
	Cin=> Carry( 	773	),
	Cout=> Carry( 	774	),
	S=> E(	761	));
			
 U775	: Somador_Exato_1 PORT MAP(
	A=> C(	839	),
	B=> E(	700	),
	Cin=> Carry( 	774	),
	Cout=> Carry( 	775	),
	S=> E(	762	));
			
 U776	: Somador_Exato_1 PORT MAP(
	A=> C(	840	),
	B=> E(	701	),
	Cin=> Carry( 	775	),
	Cout=> Carry( 	776	),
	S=> E(	763	));
			
 U777	: Somador_Exato_1 PORT MAP(
	A=> C(	841	),
	B=> E(	702	),
	Cin=> Carry( 	776	),
	Cout=> Carry( 	777	),
	S=> E(	764	));
			
 U778	: Somador_Exato_1 PORT MAP(
	A=> C(	842	),
	B=> E(	703	),
	Cin=> Carry( 	777	),
	Cout=> Carry( 	778	),
	S=> E(	765	));
			
 U779	: Somador_Exato_1 PORT MAP(
	A=> C(	843	),
	B=> E(	704	),
	Cin=> Carry( 	778	),
	Cout=> Carry( 	779	),
	S=> E(	766	));
			
 U780	: Somador_Exato_1 PORT MAP(
	A=> C(	844	),
	B=> E(	705	),
	Cin=> Carry( 	779	),
	Cout=> Carry( 	780	),
	S=> E(	767	));
			
 U781	: Somador_Exato_1 PORT MAP(
	A=> C(	845	),
	B=> E(	706	),
	Cin=> Carry( 	780	),
	Cout=> Carry( 	781	),
	S=> E(	768	));
			
 U782	: Somador_Exato_1 PORT MAP(
	A=> C(	846	),
	B=> E(	707	),
	Cin=> Carry( 	781	),
	Cout=> Carry( 	782	),
	S=> E(	769	));
			
 U783	: Somador_Exato_1 PORT MAP(
	A=> C(	847	),
	B=> E(	708	),
	Cin=> Carry( 	782	),
	Cout=> Carry( 	783	),
	S=> E(	770	));
			
 U784	: Somador_Exato_1 PORT MAP(
	A=> C(	848	),
	B=> E(	709	),
	Cin=> Carry( 	783	),
	Cout=> Carry( 	784	),
	S=> E(	771	));
			
 U785	: Somador_Exato_1 PORT MAP(
	A=> C(	849	),
	B=> E(	710	),
	Cin=> Carry( 	784	),
	Cout=> Carry( 	785	),
	S=> E(	772	));
			
 U786	: Somador_Exato_1 PORT MAP(
	A=> C(	850	),
	B=> E(	711	),
	Cin=> Carry( 	785	),
	Cout=> Carry( 	786	),
	S=> E(	773	));
			
 U787	: Somador_Exato_1 PORT MAP(
	A=> C(	851	),
	B=> E(	712	),
	Cin=> Carry( 	786	),
	Cout=> Carry( 	787	),
	S=> E(	774	));
			
 U788	: Somador_Exato_1 PORT MAP(
	A=> C(	852	),
	B=> E(	713	),
	Cin=> Carry( 	787	),
	Cout=> Carry( 	788	),
	S=> E(	775	));
			
 U789	: Somador_Exato_1 PORT MAP(
	A=> C(	853	),
	B=> E(	714	),
	Cin=> Carry( 	788	),
	Cout=> Carry( 	789	),
	S=> E(	776	));
			
 U790	: Somador_Exato_1 PORT MAP(
	A=> C(	854	),
	B=> E(	715	),
	Cin=> Carry( 	789	),
	Cout=> Carry( 	790	),
	S=> E(	777	));
			
 U791	: Somador_Exato_1 PORT MAP(
	A=> C(	855	),
	B=> E(	716	),
	Cin=> Carry( 	790	),
	Cout=> Carry( 	791	),
	S=> E(	778	));
			
 U792	: Somador_Exato_1 PORT MAP(
	A=> C(	856	),
	B=> E(	717	),
	Cin=> Carry( 	791	),
	Cout=> Carry( 	792	),
	S=> E(	779	));
			
 U793	: Somador_Exato_1 PORT MAP(
	A=> C(	857	),
	B=> E(	718	),
	Cin=> Carry( 	792	),
	Cout=> Carry( 	793	),
	S=> E(	780	));
			
 U794	: Somador_Exato_1 PORT MAP(
	A=> C(	858	),
	B=> E(	719	),
	Cin=> Carry( 	793	),
	Cout=> Carry( 	794	),
	S=> E(	781	));
			
 U795	: Somador_Exato_1 PORT MAP(
	A=> C(	859	),
	B=> E(	720	),
	Cin=> Carry( 	794	),
	Cout=> Carry( 	795	),
	S=> E(	782	));
			
 U796	: Somador_Exato_1 PORT MAP(
	A=> C(	860	),
	B=> E(	721	),
	Cin=> Carry( 	795	),
	Cout=> Carry( 	796	),
	S=> E(	783	));
			
 U797	: Somador_Exato_1 PORT MAP(
	A=> C(	861	),
	B=> E(	722	),
	Cin=> Carry( 	796	),
	Cout=> Carry( 	797	),
	S=> E(	784	));
			
 U798	: Somador_Exato_1 PORT MAP(
	A=> C(	862	),
	B=> E(	723	),
	Cin=> Carry( 	797	),
	Cout=> Carry( 	798	),
	S=> E(	785	));
			
 U799	: Somador_Exato_1 PORT MAP(
	A=> C(	863	),
	B=> E(	724	),
	Cin=> Carry( 	798	),
	Cout=> Carry( 	799	),
	S=> E(	786	));
			
 U800	: Somador_Exato_1 PORT MAP(
	A=> C(	864	),
	B=> E(	725	),
	Cin=> Carry( 	799	),
	Cout=> Carry( 	800	),
	S=> E(	787	));
			
 U801	: Somador_Exato_1 PORT MAP(
	A=> C(	865	),
	B=> E(	726	),
	Cin=> Carry( 	800	),
	Cout=> Carry( 	801	),
	S=> E(	788	));
			
 U802	: Somador_Exato_1 PORT MAP(
	A=> C(	866	),
	B=> E(	727	),
	Cin=> Carry( 	801	),
	Cout=> Carry( 	802	),
	S=> E(	789	));
			
 U803	: Somador_Exato_1 PORT MAP(
	A=> C(	867	),
	B=> E(	728	),
	Cin=> Carry( 	802	),
	Cout=> Carry( 	803	),
	S=> E(	790	));
			
 U804	: Somador_Exato_1 PORT MAP(
	A=> C(	868	),
	B=> E(	729	),
	Cin=> Carry( 	803	),
	Cout=> Carry( 	804	),
	S=> E(	791	));
			
 U805	: Somador_Exato_1 PORT MAP(
	A=> C(	869	),
	B=> E(	730	),
	Cin=> Carry( 	804	),
	Cout=> Carry( 	805	),
	S=> E(	792	));
			
 U806	: Somador_Exato_1 PORT MAP(
	A=> C(	870	),
	B=> E(	731	),
	Cin=> Carry( 	805	),
	Cout=> Carry( 	806	),
	S=> E(	793	));
			
 U807	: Somador_Exato_1 PORT MAP(
	A=> C(	871	),
	B=> E(	732	),
	Cin=> Carry( 	806	),
	Cout=> Carry( 	807	),
	S=> E(	794	));
			
 U808	: Somador_Exato_1 PORT MAP(
	A=> C(	872	),
	B=> E(	733	),
	Cin=> Carry( 	807	),
	Cout=> Carry( 	808	),
	S=> E(	795	));
			
 U809	: Somador_Exato_1 PORT MAP(
	A=> C(	873	),
	B=> E(	734	),
	Cin=> Carry( 	808	),
	Cout=> Carry( 	809	),
	S=> E(	796	));
			
 U810	: Somador_Exato_1 PORT MAP(
	A=> C(	874	),
	B=> E(	735	),
	Cin=> Carry( 	809	),
	Cout=> Carry( 	810	),
	S=> E(	797	));
			
 U811	: Somador_Exato_1 PORT MAP(
	A=> C(	875	),
	B=> E(	736	),
	Cin=> Carry( 	810	),
	Cout=> Carry( 	811	),
	S=> E(	798	));
			
 U812	: Somador_Exato_1 PORT MAP(
	A=> C(	876	),
	B=> E(	737	),
	Cin=> Carry( 	811	),
	Cout=> Carry( 	812	),
	S=> E(	799	));
			
 U813	: Somador_Exato_1 PORT MAP(
	A=> C(	877	),
	B=> E(	738	),
	Cin=> Carry( 	812	),
	Cout=> Carry( 	813	),
	S=> E(	800	));
			
 U814	: Somador_Exato_1 PORT MAP(
	A=> C(	878	),
	B=> E(	739	),
	Cin=> Carry( 	813	),
	Cout=> Carry( 	814	),
	S=> E(	801	));
			
 U815	: Somador_Exato_1 PORT MAP(
	A=> C(	879	),
	B=> E(	740	),
	Cin=> Carry( 	814	),
	Cout=> Carry( 	815	),
	S=> E(	802	));
			
 U816	: Somador_Exato_1 PORT MAP(
	A=> C(	880	),
	B=> E(	741	),
	Cin=> Carry( 	815	),
	Cout=> Carry( 	816	),
	S=> E(	803	));
			
 U817	: Somador_Exato_1 PORT MAP(
	A=> C(	881	),
	B=> E(	742	),
	Cin=> Carry( 	816	),
	Cout=> Carry( 	817	),
	S=> E(	804	));
			
 U818	: Somador_Exato_1 PORT MAP(
	A=> C(	882	),
	B=> E(	743	),
	Cin=> Carry( 	817	),
	Cout=> Carry( 	818	),
	S=> E(	805	));
			
 U819	: Somador_Exato_1 PORT MAP(
	A=> C(	883	),
	B=> E(	744	),
	Cin=> Carry( 	818	),
	Cout=> Carry( 	819	),
	S=> E(	806	));
			
 U820	: Somador_Exato_1 PORT MAP(
	A=> C(	884	),
	B=> E(	745	),
	Cin=> Carry( 	819	),
	Cout=> Carry( 	820	),
	S=> E(	807	));
			
 U821	: Somador_Exato_1 PORT MAP(
	A=> C(	885	),
	B=> E(	746	),
	Cin=> Carry( 	820	),
	Cout=> Carry( 	821	),
	S=> E(	808	));
			
 U822	: Somador_Exato_1 PORT MAP(
	A=> C(	886	),
	B=> E(	747	),
	Cin=> Carry( 	821	),
	Cout=> Carry( 	822	),
	S=> E(	809	));
			
 U823	: Somador_Exato_1 PORT MAP(
	A=> C(	887	),
	B=> E(	748	),
	Cin=> Carry( 	822	),
	Cout=> Carry( 	823	),
	S=> E(	810	));
			
 U824	: Somador_Exato_1 PORT MAP(
	A=> C(	888	),
	B=> E(	749	),
	Cin=> Carry( 	823	),
	Cout=> Carry( 	824	),
	S=> E(	811	));
			
 U825	: Somador_Exato_1 PORT MAP(
	A=> C(	889	),
	B=> E(	750	),
	Cin=> Carry( 	824	),
	Cout=> Carry( 	825	),
	S=> E(	812	));
			
 U826	: Somador_Exato_1 PORT MAP(
	A=> C(	890	),
	B=> E(	751	),
	Cin=> Carry( 	825	),
	Cout=> Carry( 	826	),
	S=> E(	813	));
			
 U827	: Somador_Exato_1 PORT MAP(
	A=> C(	891	),
	B=> E(	752	),
	Cin=> Carry( 	826	),
	Cout=> Carry( 	827	),
	S=> E(	814	));
			
 U828	: Somador_Exato_1 PORT MAP(
	A=> C(	892	),
	B=> E(	753	),
	Cin=> Carry( 	827	),
	Cout=> Carry( 	828	),
	S=> E(	815	));
			
 U829	: Somador_Exato_1 PORT MAP(
	A=> C(	893	),
	B=> E(	754	),
	Cin=> Carry( 	828	),
	Cout=> Carry( 	829	),
	S=> E(	816	));
			
 U830	: Somador_Exato_1 PORT MAP(
	A=> C(	894	),
	B=> E(	755	),
	Cin=> Carry( 	829	),
	Cout=> Carry( 	830	),
	S=> E(	817	));
			
 U831	: Somador_Exato_1 PORT MAP(
	A=> C(	895	),
	B=> Carry(	767	),
	Cin=> Carry( 	830	),
	Cout=> Carry( 	831	),
	S=> E(	818	));

			
 U832	: Somador_Exato_1 PORT MAP(
	A=> C(	896	),
	B=> E(	756	),
	Cin=> '0'	,
	Cout=> Carry( 	832	),
	S=> R(	14	));
			
 U833	: Somador_Exato_1 PORT MAP(
	A=> C(	897	),
	B=> E(	757	),
	Cin=> Carry( 	832	),
	Cout=> Carry( 	833	),
	S=> E(	819	));
			
 U834	: Somador_Exato_1 PORT MAP(
	A=> C(	898	),
	B=> E(	758	),
	Cin=> Carry( 	833	),
	Cout=> Carry( 	834	),
	S=> E(	820	));
			
 U835	: Somador_Exato_1 PORT MAP(
	A=> C(	899	),
	B=> E(	759	),
	Cin=> Carry( 	834	),
	Cout=> Carry( 	835	),
	S=> E(	821	));
			
 U836	: Somador_Exato_1 PORT MAP(
	A=> C(	900	),
	B=> E(	760	),
	Cin=> Carry( 	835	),
	Cout=> Carry( 	836	),
	S=> E(	822	));
			
 U837	: Somador_Exato_1 PORT MAP(
	A=> C(	901	),
	B=> E(	761	),
	Cin=> Carry( 	836	),
	Cout=> Carry( 	837	),
	S=> E(	823	));
			
 U838	: Somador_Exato_1 PORT MAP(
	A=> C(	902	),
	B=> E(	762	),
	Cin=> Carry( 	837	),
	Cout=> Carry( 	838	),
	S=> E(	824	));
			
 U839	: Somador_Exato_1 PORT MAP(
	A=> C(	903	),
	B=> E(	763	),
	Cin=> Carry( 	838	),
	Cout=> Carry( 	839	),
	S=> E(	825	));
			
 U840	: Somador_Exato_1 PORT MAP(
	A=> C(	904	),
	B=> E(	764	),
	Cin=> Carry( 	839	),
	Cout=> Carry( 	840	),
	S=> E(	826	));
			
 U841	: Somador_Exato_1 PORT MAP(
	A=> C(	905	),
	B=> E(	765	),
	Cin=> Carry( 	840	),
	Cout=> Carry( 	841	),
	S=> E(	827	));
			
 U842	: Somador_Exato_1 PORT MAP(
	A=> C(	906	),
	B=> E(	766	),
	Cin=> Carry( 	841	),
	Cout=> Carry( 	842	),
	S=> E(	828	));
			
 U843	: Somador_Exato_1 PORT MAP(
	A=> C(	907	),
	B=> E(	767	),
	Cin=> Carry( 	842	),
	Cout=> Carry( 	843	),
	S=> E(	829	));
			
 U844	: Somador_Exato_1 PORT MAP(
	A=> C(	908	),
	B=> E(	768	),
	Cin=> Carry( 	843	),
	Cout=> Carry( 	844	),
	S=> E(	830	));
			
 U845	: Somador_Exato_1 PORT MAP(
	A=> C(	909	),
	B=> E(	769	),
	Cin=> Carry( 	844	),
	Cout=> Carry( 	845	),
	S=> E(	831	));
			
  U846	: Somador_Exato_1 PORT MAP(
	A=> C(	910	),
	B=>E(	770	),
	Cin=> Carry( 	845	),
	Cout=> Carry( 	846	),
	S=> E(	832	));
			
 U847	: Somador_Exato_1 PORT MAP(
	A=> C(	911	),
	B=> E(	771	),
	Cin=> Carry( 	846	),
	Cout=> Carry( 	847	),
	S=> E(	833	));
			
 U848	: Somador_Exato_1 PORT MAP(
	A=> C(	912	),
	B=> E(	772	),
	Cin=> Carry( 	847	),
	Cout=> Carry( 	848	),
	S=> E(	834	));
			
 U849	: Somador_Exato_1 PORT MAP(
	A=> C(	913	),
	B=> E(	773	),
	Cin=> Carry( 	848	),
	Cout=> Carry( 	849	),
	S=> E(	835	));
			
 U850	: Somador_Exato_1 PORT MAP(
	A=> C(	914	),
	B=> E(	774	),
	Cin=> Carry( 	849	),
	Cout=> Carry( 	850	),
	S=> E(	836	));
			
 U851	: Somador_Exato_1 PORT MAP(
	A=> C(	915	),
	B=> E(	775	),
	Cin=> Carry( 	850	),
	Cout=> Carry( 	851	),
	S=> E(	837	));
			
 U852	: Somador_Exato_1 PORT MAP(
	A=> C(	916	),
	B=> E(	776	),
	Cin=> Carry( 	851	),
	Cout=> Carry( 	852	),
	S=> E(	838	));
			
 U853	: Somador_Exato_1 PORT MAP(
	A=> C(	917	),
	B=> E(	777	),
	Cin=> Carry( 	852	),
	Cout=> Carry( 	853	),
	S=> E(	839	));
			
 U854	: Somador_Exato_1 PORT MAP(
	A=> C(	918	),
	B=> E(	778	),
	Cin=> Carry( 	853	),
	Cout=> Carry( 	854	),
	S=> E(	840	));
			
 U855	: Somador_Exato_1 PORT MAP(
	A=> C(	919	),
	B=> E(	779	),
	Cin=> Carry( 	854	),
	Cout=> Carry( 	855	),
	S=> E(	841	));
			
 U856	: Somador_Exato_1 PORT MAP(
	A=> C(	920	),
	B=> E(	780	),
	Cin=> Carry( 	855	),
	Cout=> Carry( 	856	),
	S=> E(	842	));
			
 U857	: Somador_Exato_1 PORT MAP(
	A=> C(	921	),
	B=> E(	781	),
	Cin=> Carry( 	856	),
	Cout=> Carry( 	857	),
	S=> E(	843	));
			
 U858	: Somador_Exato_1 PORT MAP(
	A=> C(	922	),
	B=> E(	782	),
	Cin=> Carry( 	857	),
	Cout=> Carry( 	858	),
	S=> E(	844	));
			
 U859	: Somador_Exato_1 PORT MAP(
	A=> C(	923	),
	B=> E(	783	),
	Cin=> Carry( 	858	),
	Cout=> Carry( 	859	),
	S=> E(	845	));
			
 U860	: Somador_Exato_1 PORT MAP(
	A=> C(	924	),
	B=> E(	784	),
	Cin=> Carry( 	859	),
	Cout=> Carry( 	860	),
	S=> E(	846	));
			
 U861	: Somador_Exato_1 PORT MAP(
	A=> C(	925	),
	B=> E(	785	),
	Cin=> Carry( 	860	),
	Cout=> Carry( 	861	),
	S=> E(	847	));
			
  U862	: Somador_Exato_1 PORT MAP(
	A=> C(	926	),
	B=> E(	786	),
	Cin=> Carry( 	861	),
	Cout=> Carry( 	862	),
	S=> E(	848	));
			
 U863	: Somador_Exato_1 PORT MAP(
	A=> C(	927	),
	B=> E(	787	),
	Cin=> Carry( 	862	),
	Cout=> Carry( 	863	),
	S=> E(	849	));
			
 U864	: Somador_Exato_1 PORT MAP(
	A=> C(	928	),
	B=> E(	788	),
	Cin=> Carry( 	863	),
	Cout=> Carry( 	864	),
	S=> E(	850	));
			
 U865	: Somador_Exato_1 PORT MAP(
	A=> C(	929	),
	B=> E(	789	),
	Cin=> Carry( 	864	),
	Cout=> Carry( 	865	),
	S=> E(	851	));
			
 U866	: Somador_Exato_1 PORT MAP(
	A=> C(	930	),
	B=> E(	790	),
	Cin=> Carry( 	865	),
	Cout=> Carry( 	866	),
	S=> E(	852	));
			
 U867	: Somador_Exato_1 PORT MAP(
	A=> C(	931	),
	B=> E(	791	),
	Cin=> Carry( 	866	),
	Cout=> Carry( 	867	),
	S=> E(	853	));
			
 U868	: Somador_Exato_1 PORT MAP(
	A=> C(	932	),
	B=> E(	792	),
	Cin=> Carry( 	867	),
	Cout=> Carry( 	868	),
	S=> E(	854	));
			
 U869	: Somador_Exato_1 PORT MAP(
	A=> C(	933	),
	B=> E(	793	),
	Cin=> Carry( 	868	),
	Cout=> Carry( 	869	),
	S=> E(	855	));
			
 U870	: Somador_Exato_1 PORT MAP(
	A=> C(	934	),
	B=> E(	794	),
	Cin=> Carry( 	869	),
	Cout=> Carry( 	870	),
	S=> E(	856	));
			
 U871	: Somador_Exato_1 PORT MAP(
	A=> C(	935	),
	B=> E(	795	),
	Cin=> Carry( 	870	),
	Cout=> Carry( 	871	),
	S=> E(	857	));
			
 U872	: Somador_Exato_1 PORT MAP(
	A=> C(	936	),
	B=> E(	796	),
	Cin=> Carry( 	871	),
	Cout=> Carry( 	872	),
	S=> E(	858	));
			
 U873	: Somador_Exato_1 PORT MAP(
	A=> C(	937	),
	B=> E(	797	),
	Cin=> Carry( 	872	),
	Cout=> Carry( 	873	),
	S=> E(	859	));
			
 U874	: Somador_Exato_1 PORT MAP(
	A=> C(	938	),
	B=> E(	798	),
	Cin=> Carry( 	873	),
	Cout=> Carry( 	874	),
	S=> E(	860	));
			
 U875	: Somador_Exato_1 PORT MAP(
	A=> C(	939	),
	B=> E(	799	),
	Cin=> Carry( 	874	),
	Cout=> Carry( 	875	),
	S=> E(	861	));
			
 U876	: Somador_Exato_1 PORT MAP(
	A=> C(	940	),
	B=> E(	800	),
	Cin=> Carry( 	875	),
	Cout=> Carry( 	876	),
	S=> E(	862	));
			
 U877	: Somador_Exato_1 PORT MAP(
	A=> C(	941	),
	B=> E(	801	),
	Cin=> Carry( 	876	),
	Cout=> Carry( 	877	),
	S=> E(	863	));
			
 U878	: Somador_Exato_1 PORT MAP(
	A=> C(	942	),
	B=> E(	802	),
	Cin=> Carry( 	877	),
	Cout=> Carry( 	878	),
	S=> E(	864	));
			
 U879	: Somador_Exato_1 PORT MAP(
	A=> C(	943	),
	B=> E(	803	),
	Cin=> Carry( 	878	),
	Cout=> Carry( 	879	),
	S=> E(	865	));
			
 U880	: Somador_Exato_1 PORT MAP(
	A=> C(	944	),
	B=> E(	804	),
	Cin=> Carry( 	879	),
	Cout=> Carry( 	880	),
	S=> E(	866	));
			
 U881	: Somador_Exato_1 PORT MAP(
	A=> C(	945	),
	B=> E(	805	),
	Cin=> Carry( 	880	),
	Cout=> Carry( 	881	),
	S=> E(	867	));
			
 U882	: Somador_Exato_1 PORT MAP(
	A=> C(	946	),
	B=> E(	806	),
	Cin=> Carry( 	881	),
	Cout=> Carry( 	882	),
	S=> E(	868	));
			
 U883	: Somador_Exato_1 PORT MAP(
	A=> C(	947	),
	B=> E(	807	),
	Cin=> Carry( 	882	),
	Cout=> Carry( 	883	),
	S=> E(	869	));
			
 U884	: Somador_Exato_1 PORT MAP(
	A=> C(	948	),
	B=> E(	808	),
	Cin=> Carry( 	883	),
	Cout=> Carry( 	884	),
	S=> E(	870	));
			
 U885	: Somador_Exato_1 PORT MAP(
	A=> C(	949	),
	B=> E(	809	),
	Cin=> Carry( 	884	),
	Cout=> Carry( 	885	),
	S=> E(	871	));
			
 U886	: Somador_Exato_1 PORT MAP(
	A=> C(	950	),
	B=> E(	810	),
	Cin=> Carry( 	885	),
	Cout=> Carry( 	886	),
	S=> E(	872	));
			
 U887	: Somador_Exato_1 PORT MAP(
	A=> C(	951	),
	B=> E(	811	),
	Cin=> Carry( 	886	),
	Cout=> Carry( 	887	),
	S=> E(	873	));
			
 U888	: Somador_Exato_1 PORT MAP(
	A=> C(	952	),
	B=> E(	812	),
	Cin=> Carry( 	887	),
	Cout=> Carry( 	888	),
	S=> E(	874	));
			
 U889	: Somador_Exato_1 PORT MAP(
	A=> C(	953	),
	B=> E(	813	),
	Cin=> Carry( 	888	),
	Cout=> Carry( 	889	),
	S=> E(	875	));
			
 U890	: Somador_Exato_1 PORT MAP(
	A=> C(	954	),
	B=> E(	814	),
	Cin=> Carry( 	889	),
	Cout=> Carry( 	890	),
	S=> E(	876	));
			
 U891	: Somador_Exato_1 PORT MAP(
	A=> C(	955	),
	B=> E(	815	),
	Cin=> Carry( 	890	),
	Cout=> Carry( 	891	),
	S=> E(	877	));
			
 U892	: Somador_Exato_1 PORT MAP(
	A=> C(	956	),
	B=> E(	816	),
	Cin=> Carry( 	891	),
	Cout=> Carry( 	892	),
	S=> E(	878	));
			
 U893	: Somador_Exato_1 PORT MAP(
	A=> C(	957	),
	B=> E(	817	),
	Cin=> Carry( 	892	),
	Cout=> Carry( 	893	),
	S=> E(	879	));
			
 U894	: Somador_Exato_1 PORT MAP(
	A=> C(	958	),
	B=> E(	818	),
	Cin=> Carry( 	893	),
	Cout=> Carry( 	894	),
	S=> E(	880	));
			
 U895	: Somador_Exato_1 PORT MAP(
	A=> C(	959	),
	B=> Carry(	831	),
	Cin=> Carry( 	894	),
	Cout=> Carry( 	895	),
	S=> E(	881	));

			
 U896	: Somador_Exato_1 PORT MAP(
	A=> C(	960	),
	B=> E(	819	),
	Cin=> '0'	,
	Cout=> Carry( 	896	),
	S=> R(	15	));
			
 U897	: Somador_Exato_1 PORT MAP(
	A=> C(	961	),
	B=> E(	820	),
	Cin=> Carry( 	896	),
	Cout=> Carry( 	897	),
	S=> E(	882	));
			
 U898	: Somador_Exato_1 PORT MAP(
	A=> C(	962	),
	B=> E(	821	),
	Cin=> Carry( 	897	),
	Cout=> Carry( 	898	),
	S=> E(	883	));
			
 U899	: Somador_Exato_1 PORT MAP(
	A=> C(	963	),
	B=> E(	822	),
	Cin=> Carry( 	898	),
	Cout=> Carry( 	899	),
	S=> E(	884	));
			
 U900	: Somador_Exato_1 PORT MAP(
	A=> C(	964	),
	B=> E(	823	),
	Cin=> Carry( 	899	),
	Cout=> Carry( 	900	),
	S=> E(	885	));
			
 U901	: Somador_Exato_1 PORT MAP(
	A=> C(	965	),
	B=> E(	824	),
	Cin=> Carry( 	900	),
	Cout=> Carry( 	901	),
	S=> E(	886	));
			
 U902	: Somador_Exato_1 PORT MAP(
	A=> C(	966	),
	B=> E(	825	),
	Cin=> Carry( 	901	),
	Cout=> Carry( 	902	),
	S=> E(	887	));
			
 U903	: Somador_Exato_1 PORT MAP(
	A=> C(	967	),
	B=> E(	826	),
	Cin=> Carry( 	902	),
	Cout=> Carry( 	903	),
	S=> E(	888	));
			
 U904	: Somador_Exato_1 PORT MAP(
	A=> C(	968	),
	B=> E(	827	),
	Cin=> Carry( 	903	),
	Cout=> Carry( 	904	),
	S=> E(	889	));
			
 U905	: Somador_Exato_1 PORT MAP(
	A=> C(	969	),
	B=> E(	828	),
	Cin=> Carry( 	904	),
	Cout=> Carry( 	905	),
	S=> E(	890	));
			
 U906	: Somador_Exato_1 PORT MAP(
	A=> C(	970	),
	B=> E(	829	),
	Cin=> Carry( 	905	),
	Cout=> Carry( 	906	),
	S=> E(	891	));
			
 U907	: Somador_Exato_1 PORT MAP(
	A=> C(	971	),
	B=> E(	830	),
	Cin=> Carry( 	906	),
	Cout=> Carry( 	907	),
	S=> E(	892	));
			
 U908	: Somador_Exato_1 PORT MAP(
	A=> C(	972	),
	B=> E(	831	),
	Cin=> Carry( 	907	),
	Cout=> Carry( 	908	),
	S=> E(	893	));
			
 U909	: Somador_Exato_1 PORT MAP(
	A=> C(	973	),
	B=> E(	832	),
	Cin=> Carry( 	908	),
	Cout=> Carry( 	909	),
	S=> E(	894	));
			
 U910	: Somador_Exato_1 PORT MAP(
	A=> C(	974	),
	B=> E(	833	),
	Cin=> Carry( 	909	),
	Cout=> Carry( 	910	),
	S=> E(	895	));
			
 U911	: Somador_Exato_1 PORT MAP(
	A=> C(	975	),
	B=> E(	834	),
	Cin=> Carry( 	910	),
	Cout=> Carry( 	911	),
	S=> E(	896	));
			
 U912	: Somador_Exato_1 PORT MAP(
	A=> C(	976	),
	B=> E(	835	),
	Cin=> Carry( 	911	),
	Cout=> Carry( 	912	),
	S=> E(	897	));
			
 U913	: Somador_Exato_1 PORT MAP(
	A=> C(	977	),
	B=> E(	836	),
	Cin=> Carry( 	912	),
	Cout=> Carry( 	913	),
	S=> E(	898	));
			
 U914	: Somador_Exato_1 PORT MAP(
	A=> C(	978	),
	B=> E(	837	),
	Cin=> Carry( 	913	),
	Cout=> Carry( 	914	),
	S=> E(	899	));
			
 U915	: Somador_Exato_1 PORT MAP(
	A=> C(	979	),
	B=> E(	838	),
	Cin=> Carry( 	914	),
	Cout=> Carry( 	915	),
	S=> E(	900	));
			
 U916	: Somador_Exato_1 PORT MAP(
	A=> C(	980	),
	B=> E(	839	),
	Cin=> Carry( 	915	),
	Cout=> Carry( 	916	),
	S=> E(	901	));
			
 U917	: Somador_Exato_1 PORT MAP(
	A=> C(	981	),
	B=> E(	840	),
	Cin=> Carry( 	916	),
	Cout=> Carry( 	917	),
	S=> E(	902	));
			
 U918	: Somador_Exato_1 PORT MAP(
	A=> C(	982	),
	B=> E(	841	),
	Cin=> Carry( 	917	),
	Cout=> Carry( 	918	),
	S=> E(	903	));
			
 U919	: Somador_Exato_1 PORT MAP(
	A=> C(	983	),
	B=> E(	842	),
	Cin=> Carry( 	918	),
	Cout=> Carry( 	919	),
	S=> E(	904	));
			
 U920	: Somador_Exato_1 PORT MAP(
	A=> C(	984	),
	B=> E(	843	),
	Cin=> Carry( 	919	),
	Cout=> Carry( 	920	),
	S=> E(	905	));
			
 U921	: Somador_Exato_1 PORT MAP(
	A=> C(	985	),
	B=> E(	844	),
	Cin=> Carry( 	920	),
	Cout=> Carry( 	921	),
	S=> E(	906	));
			
 U922	: Somador_Exato_1 PORT MAP(
	A=> C(	986	),
	B=> E(	845	),
	Cin=> Carry( 	921	),
	Cout=> Carry( 	922	),
	S=> E(	907	));
			
 U923	: Somador_Exato_1 PORT MAP(
	A=> C(	987	),
	B=> E(	846	),
	Cin=> Carry( 	922	),
	Cout=> Carry( 	923	),
	S=> E(	908	));
			
 U924	: Somador_Exato_1 PORT MAP(
	A=> C(	988	),
	B=> E(	847	),
	Cin=> Carry( 	923	),
	Cout=> Carry( 	924	),
	S=> E(	909	));
			
 U925	: Somador_Exato_1 PORT MAP(
	A=> C(	989	),
	B=> E(	848	),
	Cin=> Carry( 	924	),
	Cout=> Carry( 	925	),
	S=> E(	910	));
			
 U926	: Somador_Exato_1 PORT MAP(
	A=> C(	990	),
	B=> E(	849	),
	Cin=> Carry( 	925	),
	Cout=> Carry( 	926	),
	S=> E(	911	));
			
 U927	: Somador_Exato_1 PORT MAP(
	A=> C(	991	),
	B=> E(	850	),
	Cin=> Carry( 	926	),
	Cout=> Carry( 	927	),
	S=> E(	912	));
			
 U928	: Somador_Exato_1 PORT MAP(
	A=> C(	992	),
	B=> E(	851	),
	Cin=> Carry( 	927	),
	Cout=> Carry( 	928	),
	S=> E(	913	));
			
 U929	: Somador_Exato_1 PORT MAP(
	A=> C(	993	),
	B=>E(	852	),
	Cin=> Carry( 	928	),
	Cout=> Carry( 	929	),
	S=> E(	914	));
			
 U930	: Somador_Exato_1 PORT MAP(
	A=> C(	994	),
	B=>E(	853	),
	Cin=> Carry( 	929	),
	Cout=> Carry( 	930	),
	S=> E(	915	));
			
 U931	: Somador_Exato_1 PORT MAP(
	A=> C(	995	),
	B=>E(	854	),
	Cin=> Carry( 	930	),
	Cout=> Carry( 	931	),
	S=> E(	916	));
			
 U932	: Somador_Exato_1 PORT MAP(
	A=> C(	996	),
	B=>E(	855	),
	Cin=> Carry( 	931	),
	Cout=> Carry( 	932	),
	S=> E(	917	));
			
 U933	: Somador_Exato_1 PORT MAP(
	A=> C(	997	),
	B=>E(	856	),
	Cin=> Carry( 	932	),
	Cout=> Carry( 	933	),
	S=> E(	918	));
			
 U934	: Somador_Exato_1 PORT MAP(
	A=> C(	998	),
	B=>E(	857	),
	Cin=> Carry( 	933	),
	Cout=> Carry( 	934	),
	S=> E(	919	));
			
 U935	: Somador_Exato_1 PORT MAP(
	A=> C(	999	),
	B=>E(	858	),
	Cin=> Carry( 	934	),
	Cout=> Carry( 	935	),
	S=> E(	920	));
			
 U936	: Somador_Exato_1 PORT MAP(
	A=> C(	1000	),
	B=>E(	859	),
	Cin=> Carry( 	935	),
	Cout=> Carry( 	936	),
	S=> E(	921	));
			
 U937	: Somador_Exato_1 PORT MAP(
	A=> C(	1001	),
	B=>E(	860	),
	Cin=> Carry( 	936	),
	Cout=> Carry( 	937	),
	S=> E(	922	));
			
 U938	: Somador_Exato_1 PORT MAP(
	A=> C(	1002	),
	B=>E(	861	),
	Cin=> Carry( 	937	),
	Cout=> Carry( 	938	),
	S=> E(	923	));
			
 U939	: Somador_Exato_1 PORT MAP(
	A=> C(	1003	),
	B=>E(	862	),
	Cin=> Carry( 	938	),
	Cout=> Carry( 	939	),
	S=> E(	924	));
			
 U940	: Somador_Exato_1 PORT MAP(
	A=> C(	1004	),
	B=>E(	863	),
	Cin=> Carry( 	939	),
	Cout=> Carry( 	940	),
	S=> E(	925	));
			
 U941	: Somador_Exato_1 PORT MAP(
	A=> C(	1005	),
	B=>E(	864	),
	Cin=> Carry( 	940	),
	Cout=> Carry( 	941	),
	S=> E(	926	));
			
 U942	: Somador_Exato_1 PORT MAP(
	A=> C(	1006	),
	B=>E(	865	),
	Cin=> Carry( 	941	),
	Cout=> Carry( 	942	),
	S=> E(	927	));
			
 U943	: Somador_Exato_1 PORT MAP(
	A=> C(	1007	),
	B=>E(	866	),
	Cin=> Carry( 	942	),
	Cout=> Carry( 	943	),
	S=> E(	928	));
			
 U944	: Somador_Exato_1 PORT MAP(
	A=> C(	1008	),
	B=>E(	867	),
	Cin=> Carry( 	943	),
	Cout=> Carry( 	944	),
	S=> E(	929	));
			
 U945	: Somador_Exato_1 PORT MAP(
	A=> C(	1009	),
	B=>E(	868	),
	Cin=> Carry( 	944	),
	Cout=> Carry( 	945	),
	S=> E(	930	));
			
 U946	: Somador_Exato_1 PORT MAP(
	A=> C(	1010	),
	B=>E(	869	),
	Cin=> Carry( 	945	),
	Cout=> Carry( 	946	),
	S=> E(	931	));
			
 U947	: Somador_Exato_1 PORT MAP(
	A=> C(	1011	),
	B=>E(	870	),
	Cin=> Carry( 	946	),
	Cout=> Carry( 	947	),
	S=> E(	932	));
			
 U948	: Somador_Exato_1 PORT MAP(
	A=> C(	1012	),
	B=>E(	871	),
	Cin=> Carry( 	947	),
	Cout=> Carry( 	948	),
	S=> E(	933	));
			
 U949	: Somador_Exato_1 PORT MAP(
	A=> C(	1013	),
	B=>E(	872	),
	Cin=> Carry( 	948	),
	Cout=> Carry( 	949	),
	S=> E(	934	));
			
 U950	: Somador_Exato_1 PORT MAP(
	A=> C(	1014	),
	B=>E(	873	),
	Cin=> Carry( 	949	),
	Cout=> Carry( 	950	),
	S=> E(	935	));
			
 U951	: Somador_Exato_1 PORT MAP(
	A=> C(	1015	),
	B=>E(	874	),
	Cin=> Carry( 	950	),
	Cout=> Carry( 	951	),
	S=> E(	936	));
			
 U952	: Somador_Exato_1 PORT MAP(
	A=> C(	1016	),
	B=>E(	875	),
	Cin=> Carry( 	951	),
	Cout=> Carry( 	952	),
	S=> E(	937	));
			
 U953	: Somador_Exato_1 PORT MAP(
	A=> C(	1017	),
	B=>E(	876	),
	Cin=> Carry( 	952	),
	Cout=> Carry( 	953	),
	S=> E(	938	));
			
 U954	: Somador_Exato_1 PORT MAP(
	A=> C(	1018	),
	B=>E(	877	),
	Cin=> Carry( 	953	),
	Cout=> Carry( 	954	),
	S=> E(	939	));
			
 U955	: Somador_Exato_1 PORT MAP(
	A=> C(	1019	),
	B=>E(	878	),
	Cin=> Carry( 	954	),
	Cout=> Carry( 	955	),
	S=> E(	940	));
			
 U956	: Somador_Exato_1 PORT MAP(
	A=> C(	1020	),
	B=>E(	879	),
	Cin=> Carry( 	955	),
	Cout=> Carry( 	956	),
	S=> E(	941	));
			
 U957	: Somador_Exato_1 PORT MAP(
	A=> C(	1021	),
	B=>E(	880	),
	Cin=> Carry( 	956	),
	Cout=> Carry( 	957	),
	S=> E(	942	));
			
 U958	: Somador_Exato_1 PORT MAP(
	A=> C(	1022	),
	B=>E(	881	),
	Cin=> Carry( 	957	),
	Cout=> Carry( 	958	),
	S=> E(	943	));
			
 U959	: Somador_Exato_1 PORT MAP(
	A=> C(	1023	),
	B=>Carry(	895	),
	Cin=> Carry( 	958	),
	Cout=> Carry( 	959	),
	S=> E(	944	));


			
 U960	: Somador_Exato_1 PORT MAP(
	A=> C(	1024	),
	B=>E(	882	),
	Cin=> '0',
	Cout=> Carry( 	960	),
	S=> R(	16	));
			
 U961	: Somador_Exato_1 PORT MAP(
	A=> C(	1025	),
	B=>E(	883	),
	Cin=> Carry( 	960	),
	Cout=> Carry( 	961	),
	S=> E(	945	));
			
 U962	: Somador_Exato_1 PORT MAP(
	A=> C(	1026	),
	B=>E(	884	),
	Cin=> Carry( 	961	),
	Cout=> Carry( 	962	),
	S=> E(	946	));
			
 U963	: Somador_Exato_1 PORT MAP(
	A=> C(	1027	),
	B=>E(	885	),
	Cin=> Carry( 	962	),
	Cout=> Carry( 	963	),
	S=> E(	947	));
			
 U964	: Somador_Exato_1 PORT MAP(
	A=> C(	1028	),
	B=>E(	886	),
	Cin=> Carry( 	963	),
	Cout=> Carry( 	964	),
	S=> E(	948	));
			
 U965	: Somador_Exato_1 PORT MAP(
	A=> C(	1029	),
	B=>E(	887	),
	Cin=> Carry( 	964	),
	Cout=> Carry( 	965	),
	S=> E(	949	));
			
 U966	: Somador_Exato_1 PORT MAP(
	A=> C(	1030	),
	B=>E(	888	),
	Cin=> Carry( 	965	),
	Cout=> Carry( 	966	),
	S=> E(	950	));
			
 U967	: Somador_Exato_1 PORT MAP(
	A=> C(	1031	),
	B=>E(	889	),
	Cin=> Carry( 	966	),
	Cout=> Carry( 	967	),
	S=> E(	951	));
			
 U968	: Somador_Exato_1 PORT MAP(
	A=> C(	1032	),
	B=>E(	890	),
	Cin=> Carry( 	967	),
	Cout=> Carry( 	968	),
	S=> E(	952	));
			
 U969	: Somador_Exato_1 PORT MAP(
	A=> C(	1033	),
	B=>E(	891	),
	Cin=> Carry( 	968	),
	Cout=> Carry( 	969	),
	S=> E(	953	));
			
 U970	: Somador_Exato_1 PORT MAP(
	A=> C(	1034	),
	B=>E(	892	),
	Cin=> Carry( 	969	),
	Cout=> Carry( 	970	),
	S=> E(	954	));
			
 U971	: Somador_Exato_1 PORT MAP(
	A=> C(	1035	),
	B=>E(	893	),
	Cin=> Carry( 	970	),
	Cout=> Carry( 	971	),
	S=> E(	955	));
			
 U972	: Somador_Exato_1 PORT MAP(
	A=> C(	1036	),
	B=>E(	894	),
	Cin=> Carry( 	971	),
	Cout=> Carry( 	972	),
	S=> E(	956	));
			
 U973	: Somador_Exato_1 PORT MAP(
	A=> C(	1037	),
	B=>E(	895	),
	Cin=> Carry( 	972	),
	Cout=> Carry( 	973	),
	S=> E(	957	));
			
 U974	: Somador_Exato_1 PORT MAP(
	A=> C(	1038	),
	B=>E(	896	),
	Cin=> Carry( 	973	),
	Cout=> Carry( 	974	),
	S=> E(	958	));
			
 U975	: Somador_Exato_1 PORT MAP(
	A=> C(	1039	),
	B=>E(	897	),
	Cin=> Carry( 	974	),
	Cout=> Carry( 	975	),
	S=> E(	959	));
			
 U976	: Somador_Exato_1 PORT MAP(
	A=> C(	1040	),
	B=>E(	898	),
	Cin=> Carry( 	975	),
	Cout=> Carry( 	976	),
	S=> E(	960	));
			
 U977	: Somador_Exato_1 PORT MAP(
	A=> C(	1041	),
	B=>E(	899	),
	Cin=> Carry( 	976	),
	Cout=> Carry( 	977	),
	S=> E(	961	));
			
 U978	: Somador_Exato_1 PORT MAP(
	A=> C(	1042	),
	B=>E(	900	),
	Cin=> Carry( 	977	),
	Cout=> Carry( 	978	),
	S=> E(	962	));
			
 U979	: Somador_Exato_1 PORT MAP(
	A=> C(	1043	),
	B=>E(	901	),
	Cin=> Carry( 	978	),
	Cout=> Carry( 	979	),
	S=> E(	963	));
			
 U980	: Somador_Exato_1 PORT MAP(
	A=> C(	1044	),
	B=>E(	902	),
	Cin=> Carry( 	979	),
	Cout=> Carry( 	980	),
	S=> E(	964	));
			
 U981	: Somador_Exato_1 PORT MAP(
	A=> C(	1045	),
	B=>E(	903	),
	Cin=> Carry( 	980	),
	Cout=> Carry( 	981	),
	S=> E(	965	));
			
 U982	: Somador_Exato_1 PORT MAP(
	A=> C(	1046	),
	B=>E(	904	),
	Cin=> Carry( 	981	),
	Cout=> Carry( 	982	),
	S=> E(	966	));
			
 U983	: Somador_Exato_1 PORT MAP(
	A=> C(	1047	),
	B=>E(	905	),
	Cin=> Carry( 	982	),
	Cout=> Carry( 	983	),
	S=> E(	967	));
			
 U984	: Somador_Exato_1 PORT MAP(
	A=> C(	1048	),
	B=>E(	906	),
	Cin=> Carry( 	983	),
	Cout=> Carry( 	984	),
	S=> E(	968	));
			
 U985	: Somador_Exato_1 PORT MAP(
	A=> C(	1049	),
	B=>E(	907	),
	Cin=> Carry( 	984	),
	Cout=> Carry( 	985	),
	S=> E(	969	));
			
 U986	: Somador_Exato_1 PORT MAP(
	A=> C(	1050	),
	B=>E(	908	),
	Cin=> Carry( 	985	),
	Cout=> Carry( 	986	),
	S=> E(	970	));
			
 U987	: Somador_Exato_1 PORT MAP(
	A=> C(	1051	),
	B=>E(	909	),
	Cin=> Carry( 	986	),
	Cout=> Carry( 	987	),
	S=> E(	971	));
			
 U988	: Somador_Exato_1 PORT MAP(
	A=> C(	1052	),
	B=>E(	910	),
	Cin=> Carry( 	987	),
	Cout=> Carry( 	988	),
	S=> E(	972	));
			
 U989	: Somador_Exato_1 PORT MAP(
	A=> C(	1053	),
	B=>E(	911	),
	Cin=> Carry( 	988	),
	Cout=> Carry( 	989	),
	S=> E(	973	));
			
 U990	: Somador_Exato_1 PORT MAP(
	A=> C(	1054	),
	B=>E(	912	),
	Cin=> Carry( 	989	),
	Cout=> Carry( 	990	),
	S=> E(	974	));
			
 U991	: Somador_Exato_1 PORT MAP(
	A=> C(	1055	),
	B=>E(	913	),
	Cin=> Carry( 	990	),
	Cout=> Carry( 	991	),
	S=> E(	975	));
			
 U992	: Somador_Exato_1 PORT MAP(
	A=> C(	1056	),
	B=>E(	914	),
	Cin=> Carry( 	991	),
	Cout=> Carry( 	992	),
	S=> E(	976	));
			
 U993	: Somador_Exato_1 PORT MAP(
	A=> C(	1057	),
	B=>E(	915	),
	Cin=> Carry( 	992	),
	Cout=> Carry( 	993	),
	S=> E(	977	));
			
 U994	: Somador_Exato_1 PORT MAP(
	A=> C(	1058	),
	B=>E(	916	),
	Cin=> Carry( 	993	),
	Cout=> Carry( 	994	),
	S=> E(	978	));
			
 U995	: Somador_Exato_1 PORT MAP(
	A=> C(	1059	),
	B=>E(	917	),
	Cin=> Carry( 	994	),
	Cout=> Carry( 	995	),
	S=> E(	979	));
			
 U996	: Somador_Exato_1 PORT MAP(
	A=> C(	1060	),
	B=>E(	918	),
	Cin=> Carry( 	995	),
	Cout=> Carry( 	996	),
	S=> E(	980	));
			
 U997	: Somador_Exato_1 PORT MAP(
	A=> C(	1061	),
	B=>E(	919	),
	Cin=> Carry( 	996	),
	Cout=> Carry( 	997	),
	S=> E(	981	));
			
 U998	: Somador_Exato_1 PORT MAP(
	A=> C(	1062	),
	B=>E(	920	),
	Cin=> Carry( 	997	),
	Cout=> Carry( 	998	),
	S=> E(	982	));
			
 U999	: Somador_Exato_1 PORT MAP(
	A=> C(	1063	),
	B=>E(	921	),
	Cin=> Carry( 	998	),
	Cout=> Carry( 	999	),
	S=> E(	983	));
			
 U1000	: Somador_Exato_1 PORT MAP(
	A=> C(	1064	),
	B=>E(	922	),
	Cin=> Carry( 	999	),
	Cout=> Carry( 	1000	),
	S=> E(	984	));
			
 U1001	: Somador_Exato_1 PORT MAP(
	A=> C(	1065	),
	B=>E(	923	),
	Cin=> Carry( 	1000	),
	Cout=> Carry( 	1001	),
	S=> E(	985	));
			
 U1002	: Somador_Exato_1 PORT MAP(
	A=> C(	1066	),
	B=>E(	924	),
	Cin=> Carry( 	1001	),
	Cout=> Carry( 	1002	),
	S=> E(	986	));
			
 U1003	: Somador_Exato_1 PORT MAP(
	A=> C(	1067	),
	B=>E(	925	),
	Cin=> Carry( 	1002	),
	Cout=> Carry( 	1003	),
	S=> E(	987	));
			
 U1004	: Somador_Exato_1 PORT MAP(
	A=> C(	1068	),
	B=>E(	926	),
	Cin=> Carry( 	1003	),
	Cout=> Carry( 	1004	),
	S=> E(	988	));
			
 U1005	: Somador_Exato_1 PORT MAP(
	A=> C(	1069	),
	B=>E(	927	),
	Cin=> Carry( 	1004	),
	Cout=> Carry( 	1005	),
	S=> E(	989	));
			
 U1006	: Somador_Exato_1 PORT MAP(
	A=> C(	1070	),
	B=>E(	928	),
	Cin=> Carry( 	1005	),
	Cout=> Carry( 	1006	),
	S=> E(	990	));
			
 U1007	: Somador_Exato_1 PORT MAP(
	A=> C(	1071	),
	B=>E(	929	),
	Cin=> Carry( 	1006	),
	Cout=> Carry( 	1007	),
	S=> E(	991	));
			
 U1008	: Somador_Exato_1 PORT MAP(
	A=> C(	1072	),
	B=>E(	930	),
	Cin=> Carry( 	1007	),
	Cout=> Carry( 	1008	),
	S=> E(	992	));
			
 U1009	: Somador_Exato_1 PORT MAP(
	A=> C(	1073	),
	B=>E(	931	),
	Cin=> Carry( 	1008	),
	Cout=> Carry( 	1009	),
	S=> E(	993	));
			
 U1010	: Somador_Exato_1 PORT MAP(
	A=> C(	1074	),
	B=>E(	932	),
	Cin=> Carry( 	1009	),
	Cout=> Carry( 	1010	),
	S=> E(	994	));
			
 U1011	: Somador_Exato_1 PORT MAP(
	A=> C(	1075	),
	B=>E(	933	),
	Cin=> Carry( 	1010	),
	Cout=> Carry( 	1011	),
	S=> E(	995	));
			
 U1012	: Somador_Exato_1 PORT MAP(
	A=> C(	1076	),
	B=>E(	934	),
	Cin=> Carry( 	1011	),
	Cout=> Carry( 	1012	),
	S=> E(	996	));
			
 U1013	: Somador_Exato_1 PORT MAP(
	A=> C(	1077	),
	B=>E(	935	),
	Cin=> Carry( 	1012	),
	Cout=> Carry( 	1013	),
	S=> E(	997	));
			
 U1014	: Somador_Exato_1 PORT MAP(
	A=> C(	1078	),
	B=>E(	936	),
	Cin=> Carry( 	1013	),
	Cout=> Carry( 	1014	),
	S=> E(	998	));
			
 U1015	: Somador_Exato_1 PORT MAP(
	A=> C(	1079	),
	B=>E(	937	),
	Cin=> Carry( 	1014	),
	Cout=> Carry( 	1015	),
	S=> E(	999	));
			
 U1016	: Somador_Exato_1 PORT MAP(
	A=> C(	1080	),
	B=>E(	938	),
	Cin=> Carry( 	1015	),
	Cout=> Carry( 	1016	),
	S=> E(	1000	));
			
 U1017	: Somador_Exato_1 PORT MAP(
	A=> C(	1081	),
	B=>E(	939	),
	Cin=> Carry( 	1016	),
	Cout=> Carry( 	1017	),
	S=> E(	1001	));
			
 U1018	: Somador_Exato_1 PORT MAP(
	A=> C(	1082	),
	B=>E(	940	),
	Cin=> Carry( 	1017	),
	Cout=> Carry( 	1018	),
	S=> E(	1002	));
			
 U1019	: Somador_Exato_1 PORT MAP(
	A=> C(	1083	),
	B=>E(	941	),
	Cin=> Carry( 	1018	),
	Cout=> Carry( 	1019	),
	S=> E(	1003	));
			
 U1020	: Somador_Exato_1 PORT MAP(
	A=> C(	1084	),
	B=>E(	942	),
	Cin=> Carry( 	1019	),
	Cout=> Carry( 	1020	),
	S=> E(	1004	));
			
 U1021	: Somador_Exato_1 PORT MAP(
	A=> C(	1085	),
	B=>E(	943	),
	Cin=> Carry( 	1020	),
	Cout=> Carry( 	1021	),
	S=> E(	1005	));
			
 U1022	: Somador_Exato_1 PORT MAP(
	A=> C(	1086	),
	B=>E(	944	),
	Cin=> Carry( 	1021	),
	Cout=> Carry( 	1022	),
	S=> E(	1006	));
			
 U1023	: Somador_Exato_1 PORT MAP(
	A=> C(	1087	),
	B=>Carry(	959	),
	Cin=> Carry( 	1022	),
	Cout=> Carry( 	1023	),
	S=> E(	1007	));
-------------17
			
 U1024	: Somador_Exato_1 PORT MAP(
	A=> C(	1088	),
	B=>E(	945	),
	Cin=> '0'	,
	Cout=> Carry( 	1024	),
	S=> R(	17	));
			
 U1025	: Somador_Exato_1 PORT MAP(
	A=> C(	1089	),
	B=>E(	946	),
	Cin=> Carry( 	1024	),
	Cout=> Carry( 	1025	),
	S=> E(	1008	));
			
 U1026	: Somador_Exato_1 PORT MAP(
	A=> C(	1090	),
	B=>E(	947	),
	Cin=> Carry( 	1025	),
	Cout=> Carry( 	1026	),
	S=> E(	1009	));
			
 U1027	: Somador_Exato_1 PORT MAP(
	A=> C(	1091	),
	B=>E(	948	),
	Cin=> Carry( 	1026	),
	Cout=> Carry( 	1027	),
	S=> E(	1010	));
			
 U1028	: Somador_Exato_1 PORT MAP(
	A=> C(	1092	),
	B=>E(	949	),
	Cin=> Carry( 	1027	),
	Cout=> Carry( 	1028	),
	S=> E(	1011	));
			
 U1029	: Somador_Exato_1 PORT MAP(
	A=> C(	1093	),
	B=>E(	950	),
	Cin=> Carry( 	1028	),
	Cout=> Carry( 	1029	),
	S=> E(	1012	));
			
 U1030	: Somador_Exato_1 PORT MAP(
	A=> C(	1094	),
	B=>E(	951	),
	Cin=> Carry( 	1029	),
	Cout=> Carry( 	1030	),
	S=> E(	1013	));
			
 U1031	: Somador_Exato_1 PORT MAP(
	A=> C(	1095	),
	B=>E(	952	),
	Cin=> Carry( 	1030	),
	Cout=> Carry( 	1031	),
	S=> E(	1014	));
			
 U1032	: Somador_Exato_1 PORT MAP(
	A=> C(	1096	),
	B=>E(	953	),
	Cin=> Carry( 	1031	),
	Cout=> Carry( 	1032	),
	S=> E(	1015	));
			
 U1033	: Somador_Exato_1 PORT MAP(
	A=> C(	1097	),
	B=>E(	954	),
	Cin=> Carry( 	1032	),
	Cout=> Carry( 	1033	),
	S=> E(	1016	));
			
 U1034	: Somador_Exato_1 PORT MAP(
	A=> C(	1098	),
	B=>E(	955	),
	Cin=> Carry( 	1033	),
	Cout=> Carry( 	1034	),
	S=> E(	1017	));
			
 U1035	: Somador_Exato_1 PORT MAP(
	A=> C(	1099	),
	B=>E(	956	),
	Cin=> Carry( 	1034	),
	Cout=> Carry( 	1035	),
	S=> E(	1018	));
			
 U1036	: Somador_Exato_1 PORT MAP(
	A=> C(	1100	),
	B=>E(	957	),
	Cin=> Carry( 	1035	),
	Cout=> Carry( 	1036	),
	S=> E(	1019	));
			
 U1037	: Somador_Exato_1 PORT MAP(
	A=> C(	1101	),
	B=>E(	958	),
	Cin=> Carry( 	1036	),
	Cout=> Carry( 	1037	),
	S=> E(	1020	));
			
 U1038	: Somador_Exato_1 PORT MAP(
	A=> C(	1102	),
	B=>E(	959	),
	Cin=> Carry( 	1037	),
	Cout=> Carry( 	1038	),
	S=> E(	1021	));
			
 U1039	: Somador_Exato_1 PORT MAP(
	A=> C(	1103	),
	B=>E(	960	),
	Cin=> Carry( 	1038	),
	Cout=> Carry( 	1039	),
	S=> E(	1022	));
			
 U1040	: Somador_Exato_1 PORT MAP(
	A=> C(	1104	),
	B=>E(	961	),
	Cin=> Carry( 	1039	),
	Cout=> Carry( 	1040	),
	S=> E(	1023	));
			
 U1041	: Somador_Exato_1 PORT MAP(
	A=> C(	1105	),
	B=>E(	962	),
	Cin=> Carry( 	1040	),
	Cout=> Carry( 	1041	),
	S=> E(	1024	));
			
 U1042	: Somador_Exato_1 PORT MAP(
	A=> C(	1106	),
	B=>E(	963	),
	Cin=> Carry( 	1041	),
	Cout=> Carry( 	1042	),
	S=> E(	1025	));
			
 U1043	: Somador_Exato_1 PORT MAP(
	A=> C(	1107	),
	B=>E(	964	),
	Cin=> Carry( 	1042	),
	Cout=> Carry( 	1043	),
	S=> E(	1026	));
			
 U1044	: Somador_Exato_1 PORT MAP(
	A=> C(	1108	),
	B=>E(	965	),
	Cin=> Carry( 	1043	),
	Cout=> Carry( 	1044	),
	S=> E(	1027	));
			
 U1045	: Somador_Exato_1 PORT MAP(
	A=> C(	1109	),
	B=>E(	966	),
	Cin=> Carry( 	1044	),
	Cout=> Carry( 	1045	),
	S=> E(	1028	));
			
 U1046	: Somador_Exato_1 PORT MAP(
	A=> C(	1110	),
	B=>E(	967	),
	Cin=> Carry( 	1045	),
	Cout=> Carry( 	1046	),
	S=> E(	1029	));
			
 U1047	: Somador_Exato_1 PORT MAP(
	A=> C(	1111	),
	B=>E(	968	),
	Cin=> Carry( 	1046	),
	Cout=> Carry( 	1047	),
	S=> E(	1030	));
			
 U1048	: Somador_Exato_1 PORT MAP(
	A=> C(	1112	),
	B=>E(	969	),
	Cin=> Carry( 	1047	),
	Cout=> Carry( 	1048	),
	S=> E(	1031	));
			
 U1049	: Somador_Exato_1 PORT MAP(
	A=> C(	1113	),
	B=>E(	970	),
	Cin=> Carry( 	1048	),
	Cout=> Carry( 	1049	),
	S=> E(	1032	));
			
 U1050	: Somador_Exato_1 PORT MAP(
	A=> C(	1114	),
	B=>E(	971	),
	Cin=> Carry( 	1049	),
	Cout=> Carry( 	1050	),
	S=> E(	1033	));
			
 U1051	: Somador_Exato_1 PORT MAP(
	A=> C(	1115	),
	B=>E(	972	),
	Cin=> Carry( 	1050	),
	Cout=> Carry( 	1051	),
	S=> E(	1034	));
			
 U1052	: Somador_Exato_1 PORT MAP(
	A=> C(	1116	),
	B=>E(	973	),
	Cin=> Carry( 	1051	),
	Cout=> Carry( 	1052	),
	S=> E(	1035	));
			
 U1053	: Somador_Exato_1 PORT MAP(
	A=> C(	1117	),
	B=>E(	974	),
	Cin=> Carry( 	1052	),
	Cout=> Carry( 	1053	),
	S=> E(	1036	));
			
 U1054	: Somador_Exato_1 PORT MAP(
	A=> C(	1118	),
	B=>E(	975	),
	Cin=> Carry( 	1053	),
	Cout=> Carry( 	1054	),
	S=> E(	1037	));
			
 U1055	: Somador_Exato_1 PORT MAP(
	A=> C(	1119	),
	B=>E(	976	),
	Cin=> Carry( 	1054	),
	Cout=> Carry( 	1055	),
	S=> E(	1038	));
			
 U1056	: Somador_Exato_1 PORT MAP(
	A=> C(	1120	),
	B=>E(	977	),
	Cin=> Carry( 	1055	),
	Cout=> Carry( 	1056	),
	S=> E(	1039	));
			
 U1057	: Somador_Exato_1 PORT MAP(
	A=> C(	1121	),
	B=>E(	978	),
	Cin=> Carry( 	1056	),
	Cout=> Carry( 	1057	),
	S=> E(	1040	));
			
 U1058	: Somador_Exato_1 PORT MAP(
	A=> C(	1122	),
	B=>E(	979	),
	Cin=> Carry( 	1057	),
	Cout=> Carry( 	1058	),
	S=> E(	1041	));
			
 U1059	: Somador_Exato_1 PORT MAP(
	A=> C(	1123	),
	B=>E(	980	),
	Cin=> Carry( 	1058	),
	Cout=> Carry( 	1059	),
	S=> E(	1042	));
			
 U1060	: Somador_Exato_1 PORT MAP(
	A=> C(	1124	),
	B=>E(	981	),
	Cin=> Carry( 	1059	),
	Cout=> Carry( 	1060	),
	S=> E(	1043	));
			
 U1061	: Somador_Exato_1 PORT MAP(
	A=> C(	1125	),
	B=>E(	982	),
	Cin=> Carry( 	1060	),
	Cout=> Carry( 	1061	),
	S=> E(	1044	));
			
 U1062	: Somador_Exato_1 PORT MAP(
	A=> C(	1126	),
	B=>E(	983	),
	Cin=> Carry( 	1061	),
	Cout=> Carry( 	1062	),
	S=> E(	1045	));
			
 U1063	: Somador_Exato_1 PORT MAP(
	A=> C(	1127	),
	B=>E(	984	),
	Cin=> Carry( 	1062	),
	Cout=> Carry( 	1063	),
	S=> E(	1046	));
			
 U1064	: Somador_Exato_1 PORT MAP(
	A=> C(	1128	),
	B=>E(	985	),
	Cin=> Carry( 	1063	),
	Cout=> Carry( 	1064	),
	S=> E(	1047	));
			
 U1065	: Somador_Exato_1 PORT MAP(
	A=> C(	1129	),
	B=>E(	986	),
	Cin=> Carry( 	1064	),
	Cout=> Carry( 	1065	),
	S=> E(	1048	));
			
 U1066	: Somador_Exato_1 PORT MAP(
	A=> C(	1130	),
	B=>E(	987	),
	Cin=> Carry( 	1065	),
	Cout=> Carry( 	1066	),
	S=> E(	1049	));
			
 U1067	: Somador_Exato_1 PORT MAP(
	A=> C(	1131	),
	B=>E(	988	),
	Cin=> Carry( 	1066	),
	Cout=> Carry( 	1067	),
	S=> E(	1050	));
			
 U1068	: Somador_Exato_1 PORT MAP(
	A=> C(	1132	),
	B=>E(	989	),
	Cin=> Carry( 	1067	),
	Cout=> Carry( 	1068	),
	S=> E(	1051	));
			
 U1069	: Somador_Exato_1 PORT MAP(
	A=> C(	1133	),
	B=>E(	990	),
	Cin=> Carry( 	1068	),
	Cout=> Carry( 	1069	),
	S=> E(	1052	));
			
 U1070	: Somador_Exato_1 PORT MAP(
	A=> C(	1134	),
	B=>E(	991	),
	Cin=> Carry( 	1069	),
	Cout=> Carry( 	1070	),
	S=> E(	1053	));
			
 U1071	: Somador_Exato_1 PORT MAP(
	A=> C(	1135	),
	B=>E(	992	),
	Cin=> Carry( 	1070	),
	Cout=> Carry( 	1071	),
	S=> E(	1054	));
			
 U1072	: Somador_Exato_1 PORT MAP(
	A=> C(	1136	),
	B=>E(	993	),
	Cin=> Carry( 	1071	),
	Cout=> Carry( 	1072	),
	S=> E(	1055	));
			
 U1073	: Somador_Exato_1 PORT MAP(
	A=> C(	1137	),
	B=>E(	994	),
	Cin=> Carry( 	1072	),
	Cout=> Carry( 	1073	),
	S=> E(	1056	));
			
 U1074	: Somador_Exato_1 PORT MAP(
	A=> C(	1138	),
	B=>E(	995	),
	Cin=> Carry( 	1073	),
	Cout=> Carry( 	1074	),
	S=> E(	1057	));
			
 U1075	: Somador_Exato_1 PORT MAP(
	A=> C(	1139	),
	B=>E(	996	),
	Cin=> Carry( 	1074	),
	Cout=> Carry( 	1075	),
	S=> E(	1058	));
			
 U1076	: Somador_Exato_1 PORT MAP(
	A=> C(	1140	),
	B=>E(	997	),
	Cin=> Carry( 	1075	),
	Cout=> Carry( 	1076	),
	S=> E(	1059	));
			
 U1077	: Somador_Exato_1 PORT MAP(
	A=> C(	1141	),
	B=>E(	998	),
	Cin=> Carry( 	1076	),
	Cout=> Carry( 	1077	),
	S=> E(	1060	));
			
 U1078	: Somador_Exato_1 PORT MAP(
	A=> C(	1142	),
	B=>E(	999	),
	Cin=> Carry( 	1077	),
	Cout=> Carry( 	1078	),
	S=> E(	1061	));
			
 U1079	: Somador_Exato_1 PORT MAP(
	A=> C(	1143	),
	B=>E(	1000	),
	Cin=> Carry( 	1078	),
	Cout=> Carry( 	1079	),
	S=> E(	1062	));
			
 U1080	: Somador_Exato_1 PORT MAP(
	A=> C(	1144	),
	B=>E(	1001	),
	Cin=> Carry( 	1079	),
	Cout=> Carry( 	1080	),
	S=> E(	1063	));
			
 U1081	: Somador_Exato_1 PORT MAP(
	A=> C(	1145	),
	B=>E(	1002	),
	Cin=> Carry( 	1080	),
	Cout=> Carry( 	1081	),
	S=> E(	1064	));
			
 U1082	: Somador_Exato_1 PORT MAP(
	A=> C(	1146	),
	B=>E(	1003	),
	Cin=> Carry( 	1081	),
	Cout=> Carry( 	1082	),
	S=> E(	1065	));
			
 U1083	: Somador_Exato_1 PORT MAP(
	A=> C(	1147	),
	B=>E(	1004	),
	Cin=> Carry( 	1082	),
	Cout=> Carry( 	1083	),
	S=> E(	1066	));
			
 U1084	: Somador_Exato_1 PORT MAP(
	A=> C(	1148	),
	B=>E(	1005	),
	Cin=> Carry( 	1083	),
	Cout=> Carry( 	1084	),
	S=> E(	1067	));
			
 U1085	: Somador_Exato_1 PORT MAP(
	A=> C(	1149	),
	B=>E(	1006	),
	Cin=> Carry( 	1084	),
	Cout=> Carry( 	1085	),
	S=> E(	1068	));
			
 U1086	: Somador_Exato_1 PORT MAP(
	A=> C(	1150	),
	B=>E(	1007	),
	Cin=> Carry( 	1085	),
	Cout=> Carry( 	1086	),
	S=> E(	1069	));
			
 U1087	: Somador_Exato_1 PORT MAP(
	A=> C(	1151	),
	B=>Carry(	1023	),
	Cin=> Carry( 	1086	),
	Cout=> Carry( 	1087	),
	S=> E(	1070	));
-----------------
	
			
 U1088	: Somador_Exato_1 PORT MAP(
	A=> C(	1152	),
	B=>E(	1008	),
	Cin=> '0'	,
	Cout=> Carry( 	1088	),
	S=> R(	18	));
			
 U1089	: Somador_Exato_1 PORT MAP(
	A=> C(	1153	),
	B=>E(	1009	),
	Cin=> Carry( 	1088	),
	Cout=> Carry( 	1089	),
	S=> E(	1071	));
			
 U1090	: Somador_Exato_1 PORT MAP(
	A=> C(	1154	),
	B=>E(	1010	),
	Cin=> Carry( 	1089	),
	Cout=> Carry( 	1090	),
	S=> E(	1072	));
			
 U1091	: Somador_Exato_1 PORT MAP(
	A=> C(	1155	),
	B=>E(	1011	),
	Cin=> Carry( 	1090	),
	Cout=> Carry( 	1091	),
	S=> E(	1073	));
			
 U1092	: Somador_Exato_1 PORT MAP(
	A=> C(	1156	),
	B=>E(	1012	),
	Cin=> Carry( 	1091	),
	Cout=> Carry( 	1092	),
	S=> E(	1074	));
			
 U1093	: Somador_Exato_1 PORT MAP(
	A=> C(	1157	),
	B=>E(	1013	),
	Cin=> Carry( 	1092	),
	Cout=> Carry( 	1093	),
	S=> E(	1075	));
			
 U1094	: Somador_Exato_1 PORT MAP(
	A=> C(	1158	),
	B=>E(	1014	),
	Cin=> Carry( 	1093	),
	Cout=> Carry( 	1094	),
	S=> E(	1076	));
			
 U1095	: Somador_Exato_1 PORT MAP(
	A=> C(	1159	),
	B=>E(	1015	),
	Cin=> Carry( 	1094	),
	Cout=> Carry( 	1095	),
	S=> E(	1077	));
			
 U1096	: Somador_Exato_1 PORT MAP(
	A=> C(	1160	),
	B=>E(	1016	),
	Cin=> Carry( 	1095	),
	Cout=> Carry( 	1096	),
	S=> E(	1078	));
			
 U1097	: Somador_Exato_1 PORT MAP(
	A=> C(	1161	),
	B=>E(	1017	),
	Cin=> Carry( 	1096	),
	Cout=> Carry( 	1097	),
	S=> E(	1079	));
			
 U1098	: Somador_Exato_1 PORT MAP(
	A=> C(	1162	),
	B=>E(	1018	),
	Cin=> Carry( 	1097	),
	Cout=> Carry( 	1098	),
	S=> E(	1080	));
			
 U1099	: Somador_Exato_1 PORT MAP(
	A=> C(	1163	),
	B=>E(	1019	),
	Cin=> Carry( 	1098	),
	Cout=> Carry( 	1099	),
	S=> E(	1081	));
			
 U1100	: Somador_Exato_1 PORT MAP(
	A=> C(	1164	),
	B=>E(	1020	),
	Cin=> Carry( 	1099	),
	Cout=> Carry( 	1100	),
	S=> E(	1082	));
			
 U1101	: Somador_Exato_1 PORT MAP(
	A=> C(	1165	),
	B=>E(	1021	),
	Cin=> Carry( 	1100	),
	Cout=> Carry( 	1101	),
	S=> E(	1083	));
			
 U1102	: Somador_Exato_1 PORT MAP(
	A=> C(	1166	),
	B=>E(	1022	),
	Cin=> Carry( 	1101	),
	Cout=> Carry( 	1102	),
	S=> E(	1084	));
			
 U1103	: Somador_Exato_1 PORT MAP(
	A=> C(	1167	),
	B=>E(	1023	),
	Cin=> Carry( 	1102	),
	Cout=> Carry( 	1103	),
	S=> E(	1085	));
			
 U1104	: Somador_Exato_1 PORT MAP(
	A=> C(	1168	),
	B=>E(	1024	),
	Cin=> Carry( 	1103	),
	Cout=> Carry( 	1104	),
	S=> E(	1086	));
			
 U1105	: Somador_Exato_1 PORT MAP(
	A=> C(	1169	),
	B=>E(	1025	),
	Cin=> Carry( 	1104	),
	Cout=> Carry( 	1105	),
	S=> E(	1087	));
			
 U1106	: Somador_Exato_1 PORT MAP(
	A=> C(	1170	),
	B=>E(	1026	),
	Cin=> Carry( 	1105	),
	Cout=> Carry( 	1106	),
	S=> E(	1088	));
			
 U1107	: Somador_Exato_1 PORT MAP(
	A=> C(	1171	),
	B=>E(	1027	),
	Cin=> Carry( 	1106	),
	Cout=> Carry( 	1107	),
	S=> E(	1089	));
			
 U1108	: Somador_Exato_1 PORT MAP(
	A=> C(	1172	),
	B=>E(	1028	),
	Cin=> Carry( 	1107	),
	Cout=> Carry( 	1108	),
	S=> E(	1090	));
			
 U1109	: Somador_Exato_1 PORT MAP(
	A=> C(	1173	),
	B=>E(	1029	),
	Cin=> Carry( 	1108	),
	Cout=> Carry( 	1109	),
	S=> E(	1091	));
			
 U1110	: Somador_Exato_1 PORT MAP(
	A=> C(	1174	),
	B=>E(	1030	),
	Cin=> Carry( 	1109	),
	Cout=> Carry( 	1110	),
	S=> E(	1092	));
			
 U1111	: Somador_Exato_1 PORT MAP(
	A=> C(	1175	),
	B=>E(	1031	),
	Cin=> Carry( 	1110	),
	Cout=> Carry( 	1111	),
	S=> E(	1093	));
			
 U1112	: Somador_Exato_1 PORT MAP(
	A=> C(	1176	),
	B=>E(	1032	),
	Cin=> Carry( 	1111	),
	Cout=> Carry( 	1112	),
	S=> E(	1094	));
			
 U1113	: Somador_Exato_1 PORT MAP(
	A=> C(	1177	),
	B=>E(	1033	),
	Cin=> Carry( 	1112	),
	Cout=> Carry( 	1113	),
	S=> E(	1095	));
			
 U1114	: Somador_Exato_1 PORT MAP(
	A=> C(	1178	),
	B=>E(	1034	),
	Cin=> Carry( 	1113	),
	Cout=> Carry( 	1114	),
	S=> E(	1096	));
			
 U1115	: Somador_Exato_1 PORT MAP(
	A=> C(	1179	),
	B=>E(	1035	),
	Cin=> Carry( 	1114	),
	Cout=> Carry( 	1115	),
	S=> E(	1097	));
			
 U1116	: Somador_Exato_1 PORT MAP(
	A=> C(	1180	),
	B=>E(	1036	),
	Cin=> Carry( 	1115	),
	Cout=> Carry( 	1116	),
	S=> E(	1098	));
			
 U1117	: Somador_Exato_1 PORT MAP(
	A=> C(	1181	),
	B=>E(	1037	),
	Cin=> Carry( 	1116	),
	Cout=> Carry( 	1117	),
	S=> E(	1099	));
			
 U1118	: Somador_Exato_1 PORT MAP(
	A=> C(	1182	),
	B=>E(	1038	),
	Cin=> Carry( 	1117	),
	Cout=> Carry( 	1118	),
	S=> E(	1100	));
			
 U1119	: Somador_Exato_1 PORT MAP(
	A=> C(	1183	),
	B=>E(	1039	),
	Cin=> Carry( 	1118	),
	Cout=> Carry( 	1119	),
	S=> E(	1101	));
			
 U1120	: Somador_Exato_1 PORT MAP(
	A=> C(	1184	),
	B=>E(	1040	),
	Cin=> Carry( 	1119	),
	Cout=> Carry( 	1120	),
	S=> E(	1102	));
			
 U1121	: Somador_Exato_1 PORT MAP(
	A=> C(	1185	),
	B=>E(	1041	),
	Cin=> Carry( 	1120	),
	Cout=> Carry( 	1121	),
	S=> E(	1103	));
			
 U1122	: Somador_Exato_1 PORT MAP(
	A=> C(	1186	),
	B=>E(	1042	),
	Cin=> Carry( 	1121	),
	Cout=> Carry( 	1122	),
	S=> E(	1104	));
			
 U1123	: Somador_Exato_1 PORT MAP(
	A=> C(	1187	),
	B=>E(	1043	),
	Cin=> Carry( 	1122	),
	Cout=> Carry( 	1123	),
	S=> E(	1105	));
			
 U1124	: Somador_Exato_1 PORT MAP(
	A=> C(	1188	),
	B=>E(	1044	),
	Cin=> Carry( 	1123	),
	Cout=> Carry( 	1124	),
	S=> E(	1106	));
			
 U1125	: Somador_Exato_1 PORT MAP(
	A=> C(	1189	),
	B=>E(	1045	),
	Cin=> Carry( 	1124	),
	Cout=> Carry( 	1125	),
	S=> E(	1107	));
			
 U1126	: Somador_Exato_1 PORT MAP(
	A=> C(	1190	),
	B=>E(	1046	),
	Cin=> Carry( 	1125	),
	Cout=> Carry( 	1126	),
	S=> E(	1108	));
			
 U1127	: Somador_Exato_1 PORT MAP(
	A=> C(	1191	),
	B=>E(	1047	),
	Cin=> Carry( 	1126	),
	Cout=> Carry( 	1127	),
	S=> E(	1109	));
			
 U1128	: Somador_Exato_1 PORT MAP(
	A=> C(	1192	),
	B=>E(	1048	),
	Cin=> Carry( 	1127	),
	Cout=> Carry( 	1128	),
	S=> E(	1110	));
			
 U1129	: Somador_Exato_1 PORT MAP(
	A=> C(	1193	),
	B=>E(	1049	),
	Cin=> Carry( 	1128	),
	Cout=> Carry( 	1129	),
	S=> E(	1111	));
			
 U1130	: Somador_Exato_1 PORT MAP(
	A=> C(	1194	),
	B=>E(	1050	),
	Cin=> Carry( 	1129	),
	Cout=> Carry( 	1130	),
	S=> E(	1112	));
			
 U1131	: Somador_Exato_1 PORT MAP(
	A=> C(	1195	),
	B=>E(	1051	),
	Cin=> Carry( 	1130	),
	Cout=> Carry( 	1131	),
	S=> E(	1113	));
			
 U1132	: Somador_Exato_1 PORT MAP(
	A=> C(	1196	),
	B=>E(	1052	),
	Cin=> Carry( 	1131	),
	Cout=> Carry( 	1132	),
	S=> E(	1114	));
			
 U1133	: Somador_Exato_1 PORT MAP(
	A=> C(	1197	),
	B=>E(	1053	),
	Cin=> Carry( 	1132	),
	Cout=> Carry( 	1133	),
	S=> E(	1115	));
			
 U1134	: Somador_Exato_1 PORT MAP(
	A=> C(	1198	),
	B=>E(	1054	),
	Cin=> Carry( 	1133	),
	Cout=> Carry( 	1134	),
	S=> E(	1116	));
			
 U1135	: Somador_Exato_1 PORT MAP(
	A=> C(	1199	),
	B=>E(	1055	),
	Cin=> Carry( 	1134	),
	Cout=> Carry( 	1135	),
	S=> E(	1117	));
			
 U1136	: Somador_Exato_1 PORT MAP(
	A=> C(	1200	),
	B=>E(	1056	),
	Cin=> Carry( 	1135	),
	Cout=> Carry( 	1136	),
	S=> E(	1118	));
			
 U1137	: Somador_Exato_1 PORT MAP(
	A=> C(	1201	),
	B=>E(	1057	),
	Cin=> Carry( 	1136	),
	Cout=> Carry( 	1137	),
	S=> E(	1119	));
			
 U1138	: Somador_Exato_1 PORT MAP(
	A=> C(	1202	),
	B=>E(	1058	),
	Cin=> Carry( 	1137	),
	Cout=> Carry( 	1138	),
	S=> E(	1120	));
			
 U1139	: Somador_Exato_1 PORT MAP(
	A=> C(	1203	),
	B=>E(	1059	),
	Cin=> Carry( 	1138	),
	Cout=> Carry( 	1139	),
	S=> E(	1121	));
			
 U1140	: Somador_Exato_1 PORT MAP(
	A=> C(	1204	),
	B=>E(	1060	),
	Cin=> Carry( 	1139	),
	Cout=> Carry( 	1140	),
	S=> E(	1122	));
			
 U1141	: Somador_Exato_1 PORT MAP(
	A=> C(	1205	),
	B=>E(	1061	),
	Cin=> Carry( 	1140	),
	Cout=> Carry( 	1141	),
	S=> E(	1123	));
			
 U1142	: Somador_Exato_1 PORT MAP(
	A=> C(	1206	),
	B=>E(	1062	),
	Cin=> Carry( 	1141	),
	Cout=> Carry( 	1142	),
	S=> E(	1124	));
			
 U1143	: Somador_Exato_1 PORT MAP(
	A=> C(	1207	),
	B=>E(	1063	),
	Cin=> Carry( 	1142	),
	Cout=> Carry( 	1143	),
	S=> E(	1125	));
			
 U1144	: Somador_Exato_1 PORT MAP(
	A=> C(	1208	),
	B=>E(	1064	),
	Cin=> Carry( 	1143	),
	Cout=> Carry( 	1144	),
	S=> E(	1126	));
			
 U1145	: Somador_Exato_1 PORT MAP(
	A=> C(	1209	),
	B=>E(	1065	),
	Cin=> Carry( 	1144	),
	Cout=> Carry( 	1145	),
	S=> E(	1127	));
			
 U1146	: Somador_Exato_1 PORT MAP(
	A=> C(	1210	),
	B=>E(	1066	),
	Cin=> Carry( 	1145	),
	Cout=> Carry( 	1146	),
	S=> E(	1128	));
			
 U1147	: Somador_Exato_1 PORT MAP(
	A=> C(	1211	),
	B=>E(	1067	),
	Cin=> Carry( 	1146	),
	Cout=> Carry( 	1147	),
	S=> E(	1129	));
			
 U1148	: Somador_Exato_1 PORT MAP(
	A=> C(	1212	),
	B=>E(	1068	),
	Cin=> Carry( 	1147	),
	Cout=> Carry( 	1148	),
	S=> E(	1130	));
			
 U1149	: Somador_Exato_1 PORT MAP(
	A=> C(	1213	),
	B=>E(	1069	),
	Cin=> Carry( 	1148	),
	Cout=> Carry( 	1149	),
	S=> E(	1131	));
			
 U1150	: Somador_Exato_1 PORT MAP(
	A=> C(	1214	),
	B=>E(	1070	),
	Cin=> Carry( 	1149	),
	Cout=> Carry( 	1150	),
	S=> E(	1132	));
			
 U1151	: Somador_Exato_1 PORT MAP(
	A=> C(	1215	),
	B=>Carry(	1087	),
	Cin=> Carry( 	1150	),
	Cout=> Carry( 	1151	),
	S=> E(	1133	));

			
 U1152	: Somador_Exato_1 PORT MAP(
	A=> C(	1216	),
	B=>E(	1071	),
	Cin=> '0'	,
	Cout=> Carry( 	1152	),
	S=> R(	19	));
			
 U1153	: Somador_Exato_1 PORT MAP(
	A=> C(	1217	),
	B=>E(	1072	),
	Cin=> Carry( 	1152	),
	Cout=> Carry( 	1153	),
	S=> E(	1134	));
			
 U1154	: Somador_Exato_1 PORT MAP(
	A=> C(	1218	),
	B=>E(	1073	),
	Cin=> Carry( 	1153	),
	Cout=> Carry( 	1154	),
	S=> E(	1135	));
			
 U1155	: Somador_Exato_1 PORT MAP(
	A=> C(	1219	),
	B=>E(	1074	),
	Cin=> Carry( 	1154	),
	Cout=> Carry( 	1155	),
	S=> E(	1136	));
			
 U1156	: Somador_Exato_1 PORT MAP(
	A=> C(	1220	),
	B=>E(	1075	),
	Cin=> Carry( 	1155	),
	Cout=> Carry( 	1156	),
	S=> E(	1137	));
			
 U1157	: Somador_Exato_1 PORT MAP(
	A=> C(	1221	),
	B=>E(	1076	),
	Cin=> Carry( 	1156	),
	Cout=> Carry( 	1157	),
	S=> E(	1138	));
			
 U1158	: Somador_Exato_1 PORT MAP(
	A=> C(	1222	),
	B=>E(	1077	),
	Cin=> Carry( 	1157	),
	Cout=> Carry( 	1158	),
	S=> E(	1139	));
			
 U1159	: Somador_Exato_1 PORT MAP(
	A=> C(	1223	),
	B=>E(	1078	),
	Cin=> Carry( 	1158	),
	Cout=> Carry( 	1159	),
	S=> E(	1140	));
			
 U1160	: Somador_Exato_1 PORT MAP(
	A=> C(	1224	),
	B=>E(	1079	),
	Cin=> Carry( 	1159	),
	Cout=> Carry( 	1160	),
	S=> E(	1141	));
			
 U1161	: Somador_Exato_1 PORT MAP(
	A=> C(	1225	),
	B=>E(	1080	),
	Cin=> Carry( 	1160	),
	Cout=> Carry( 	1161	),
	S=> E(	1142	));
			
 U1162	: Somador_Exato_1 PORT MAP(
	A=> C(	1226	),
	B=>E(	1081	),
	Cin=> Carry( 	1161	),
	Cout=> Carry( 	1162	),
	S=> E(	1143	));
			
 U1163	: Somador_Exato_1 PORT MAP(
	A=> C(	1227	),
	B=>E(	1082	),
	Cin=> Carry( 	1162	),
	Cout=> Carry( 	1163	),
	S=> E(	1144	));
			
 U1164	: Somador_Exato_1 PORT MAP(
	A=> C(	1228	),
	B=>E(	1083	),
	Cin=> Carry( 	1163	),
	Cout=> Carry( 	1164	),
	S=> E(	1145	));
			
 U1165	: Somador_Exato_1 PORT MAP(
	A=> C(	1229	),
	B=>E(	1084	),
	Cin=> Carry( 	1164	),
	Cout=> Carry( 	1165	),
	S=> E(	1146	));
			
 U1166	: Somador_Exato_1 PORT MAP(
	A=> C(	1230	),
	B=>E(	1085	),
	Cin=> Carry( 	1165	),
	Cout=> Carry( 	1166	),
	S=> E(	1147	));
			
 U1167	: Somador_Exato_1 PORT MAP(
	A=> C(	1231	),
	B=>E(	1086	),
	Cin=> Carry( 	1166	),
	Cout=> Carry( 	1167	),
	S=> E(	1148	));
			
 U1168	: Somador_Exato_1 PORT MAP(
	A=> C(	1232	),
	B=>E(	1087	),
	Cin=> Carry( 	1167	),
	Cout=> Carry( 	1168	),
	S=> E(	1149	));
			
 U1169	: Somador_Exato_1 PORT MAP(
	A=> C(	1233	),
	B=>E(	1088	),
	Cin=> Carry( 	1168	),
	Cout=> Carry( 	1169	),
	S=> E(	1150	));
			
 U1170	: Somador_Exato_1 PORT MAP(
	A=> C(	1234	),
	B=>E(	1089	),
	Cin=> Carry( 	1169	),
	Cout=> Carry( 	1170	),
	S=> E(	1151	));
			
 U1171	: Somador_Exato_1 PORT MAP(
	A=> C(	1235	),
	B=>E(	1090	),
	Cin=> Carry( 	1170	),
	Cout=> Carry( 	1171	),
	S=> E(	1152	));
			
 U1172	: Somador_Exato_1 PORT MAP(
	A=> C(	1236	),
	B=>E(	1091	),
	Cin=> Carry( 	1171	),
	Cout=> Carry( 	1172	),
	S=> E(	1153	));
			
 U1173	: Somador_Exato_1 PORT MAP(
	A=> C(	1237	),
	B=>E(	1092	),
	Cin=> Carry( 	1172	),
	Cout=> Carry( 	1173	),
	S=> E(	1154	));
			
 U1174	: Somador_Exato_1 PORT MAP(
	A=> C(	1238	),
	B=>E(	1093	),
	Cin=> Carry( 	1173	),
	Cout=> Carry( 	1174	),
	S=> E(	1155	));
			
 U1175	: Somador_Exato_1 PORT MAP(
	A=> C(	1239	),
	B=>E(	1094	),
	Cin=> Carry( 	1174	),
	Cout=> Carry( 	1175	),
	S=> E(	1156	));
			
 U1176	: Somador_Exato_1 PORT MAP(
	A=> C(	1240	),
	B=>E(	1095	),
	Cin=> Carry( 	1175	),
	Cout=> Carry( 	1176	),
	S=> E(	1157	));
			
 U1177	: Somador_Exato_1 PORT MAP(
	A=> C(	1241	),
	B=>E(	1096	),
	Cin=> Carry( 	1176	),
	Cout=> Carry( 	1177	),
	S=> E(	1158	));
			
 U1178	: Somador_Exato_1 PORT MAP(
	A=> C(	1242	),
	B=>E(	1097	),
	Cin=> Carry( 	1177	),
	Cout=> Carry( 	1178	),
	S=> E(	1159	));
			
 U1179	: Somador_Exato_1 PORT MAP(
	A=> C(	1243	),
	B=>E(	1098	),
	Cin=> Carry( 	1178	),
	Cout=> Carry( 	1179	),
	S=> E(	1160	));
			
 U1180	: Somador_Exato_1 PORT MAP(
	A=> C(	1244	),
	B=>E(	1099	),
	Cin=> Carry( 	1179	),
	Cout=> Carry( 	1180	),
	S=> E(	1161	));
			
 U1181	: Somador_Exato_1 PORT MAP(
	A=> C(	1245	),
	B=>E(	1100	),
	Cin=> Carry( 	1180	),
	Cout=> Carry( 	1181	),
	S=> E(	1162	));
			
 U1182	: Somador_Exato_1 PORT MAP(
	A=> C(	1246	),
	B=>E(	1101	),
	Cin=> Carry( 	1181	),
	Cout=> Carry( 	1182	),
	S=> E(	1163	));
			
 U1183	: Somador_Exato_1 PORT MAP(
	A=> C(	1247	),
	B=>E(	1102	),
	Cin=> Carry( 	1182	),
	Cout=> Carry( 	1183	),
	S=> E(	1164	));
			
 U1184	: Somador_Exato_1 PORT MAP(
	A=> C(	1248	),
	B=>E(	1103	),
	Cin=> Carry( 	1183	),
	Cout=> Carry( 	1184	),
	S=> E(	1165	));
			
 U1185	: Somador_Exato_1 PORT MAP(
	A=> C(	1249	),
	B=>E(	1104	),
	Cin=> Carry( 	1184	),
	Cout=> Carry( 	1185	),
	S=> E(	1166	));
			
 U1186	: Somador_Exato_1 PORT MAP(
	A=> C(	1250	),
	B=>E(	1105	),
	Cin=> Carry( 	1185	),
	Cout=> Carry( 	1186	),
	S=> E(	1167	));
			
 U1187	: Somador_Exato_1 PORT MAP(
	A=> C(	1251	),
	B=>E(	1106	),
	Cin=> Carry( 	1186	),
	Cout=> Carry( 	1187	),
	S=> E(	1168	));
			
 U1188	: Somador_Exato_1 PORT MAP(
	A=> C(	1252	),
	B=>E(	1107	),
	Cin=> Carry( 	1187	),
	Cout=> Carry( 	1188	),
	S=> E(	1169	));
			
 U1189	: Somador_Exato_1 PORT MAP(
	A=> C(	1253	),
	B=>E(	1108	),
	Cin=> Carry( 	1188	),
	Cout=> Carry( 	1189	),
	S=> E(	1170	));
			
 U1190	: Somador_Exato_1 PORT MAP(
	A=> C(	1254	),
	B=>E(	1109	),
	Cin=> Carry( 	1189	),
	Cout=> Carry( 	1190	),
	S=> E(	1171	));
			
 U1191	: Somador_Exato_1 PORT MAP(
	A=> C(	1255	),
	B=>E(	1110	),
	Cin=> Carry( 	1190	),
	Cout=> Carry( 	1191	),
	S=> E(	1172	));
			
 U1192	: Somador_Exato_1 PORT MAP(
	A=> C(	1256	),
	B=>E(	1111	),
	Cin=> Carry( 	1191	),
	Cout=> Carry( 	1192	),
	S=> E(	1173	));
			
 U1193	: Somador_Exato_1 PORT MAP(
	A=> C(	1257	),
	B=>E(	1112	),
	Cin=> Carry( 	1192	),
	Cout=> Carry( 	1193	),
	S=> E(	1174	));
			
 U1194	: Somador_Exato_1 PORT MAP(
	A=> C(	1258	),
	B=>E(	1113	),
	Cin=> Carry( 	1193	),
	Cout=> Carry( 	1194	),
	S=> E(	1175	));
			
 U1195	: Somador_Exato_1 PORT MAP(
	A=> C(	1259	),
	B=>E(	1114	),
	Cin=> Carry( 	1194	),
	Cout=> Carry( 	1195	),
	S=> E(	1176	));
			
 U1196	: Somador_Exato_1 PORT MAP(
	A=> C(	1260	),
	B=>E(	1115	),
	Cin=> Carry( 	1195	),
	Cout=> Carry( 	1196	),
	S=> E(	1177	));
			
 U1197	: Somador_Exato_1 PORT MAP(
	A=> C(	1261	),
	B=>E(	1116	),
	Cin=> Carry( 	1196	),
	Cout=> Carry( 	1197	),
	S=> E(	1178	));
			
 U1198	: Somador_Exato_1 PORT MAP(
	A=> C(	1262	),
	B=>E(	1117	),
	Cin=> Carry( 	1197	),
	Cout=> Carry( 	1198	),
	S=> E(	1179	));
			
 U1199	: Somador_Exato_1 PORT MAP(
	A=> C(	1263	),
	B=>E(	1118	),
	Cin=> Carry( 	1198	),
	Cout=> Carry( 	1199	),
	S=> E(	1180	));
			
 U1200	: Somador_Exato_1 PORT MAP(
	A=> C(	1264	),
	B=>E(	1119	),
	Cin=> Carry( 	1199	),
	Cout=> Carry( 	1200	),
	S=> E(	1181	));
			
 U1201	: Somador_Exato_1 PORT MAP(
	A=> C(	1265	),
	B=>E(	1120	),
	Cin=> Carry( 	1200	),
	Cout=> Carry( 	1201	),
	S=> E(	1182	));
			
 U1202	: Somador_Exato_1 PORT MAP(
	A=> C(	1266	),
	B=>E(	1121	),
	Cin=> Carry( 	1201	),
	Cout=> Carry( 	1202	),
	S=> E(	1183	));
			
 U1203	: Somador_Exato_1 PORT MAP(
	A=> C(	1267	),
	B=>E(	1122	),
	Cin=> Carry( 	1202	),
	Cout=> Carry( 	1203	),
	S=> E(	1184	));
			
 U1204	: Somador_Exato_1 PORT MAP(
	A=> C(	1268	),
	B=>E(	1123	),
	Cin=> Carry( 	1203	),
	Cout=> Carry( 	1204	),
	S=> E(	1185	));
			
 U1205	: Somador_Exato_1 PORT MAP(
	A=> C(	1269	),
	B=>E(	1124	),
	Cin=> Carry( 	1204	),
	Cout=> Carry( 	1205	),
	S=> E(	1186	));
			
U1206	: Somador_Exato_1 PORT MAP(
	A=> C(	1270	),
	B=>E(	1125	),
	Cin=> Carry( 	1205	),
	Cout=> Carry( 	1206	),
	S=> E(	1187	));
			
 U1207	: Somador_Exato_1 PORT MAP(
	A=> C(	1271	),
	B=>E(	1126	),
	Cin=> Carry( 	1206	),
	Cout=> Carry( 	1207	),
	S=> E(	1188	));
			
 U1208	: Somador_Exato_1 PORT MAP(
	A=> C(	1272	),
	B=>E(	1127	),
	Cin=> Carry( 	1207	),
	Cout=> Carry( 	1208	),
	S=> E(	1189	));
			
 U1209	: Somador_Exato_1 PORT MAP(
	A=> C(	1273	),
	B=>E(	1128	),
	Cin=> Carry( 	1208	),
	Cout=> Carry( 	1209	),
	S=> E(	1190	));
			
 U1210	: Somador_Exato_1 PORT MAP(
	A=> C(	1274	),
	B=>E(	1129	),
	Cin=> Carry( 	1209	),
	Cout=> Carry( 	1210	),
	S=> E(	1191	));
			
 U1211	: Somador_Exato_1 PORT MAP(
	A=> C(	1275	),
	B=>E(	1130	),
	Cin=> Carry( 	1210	),
	Cout=> Carry( 	1211	),
	S=> E(	1192	));
			
 U1212	: Somador_Exato_1 PORT MAP(
	A=> C(	1276	),
	B=>E(	1131	),
	Cin=> Carry( 	1211	),
	Cout=> Carry( 	1212	),
	S=> E(	1193	));
			
 U1213	: Somador_Exato_1 PORT MAP(
	A=> C(	1277	),
	B=>E(	1132	),
	Cin=> Carry( 	1212	),
	Cout=> Carry( 	1213	),
	S=> E(	1194	));
			
 U1214	: Somador_Exato_1 PORT MAP(
	A=> C(	1278	),
	B=>E(	1133	),
	Cin=> Carry( 	1213	),
	Cout=> Carry( 	1214	),
	S=> E(	1195	));
			
 U1215	: Somador_Exato_1 PORT MAP(
	A=> C(	1279	),
	B=>Carry(	1151	),
	Cin=> Carry( 	1214	),
	Cout=> Carry( 	1215	),
	S=> E(	1196	));

			
 U1216	: Somador_Exato_1 PORT MAP(
	A=> C(	1280	),
	B=>E(	1134	),
	Cin=> '0'	,
	Cout=> Carry( 	1216	),
	S=> R(	20	));
			
 U1217	: Somador_Exato_1 PORT MAP(
	A=> C(	1281	),
	B=>E(	1135	),
	Cin=> Carry( 	1216	),
	Cout=> Carry( 	1217	),
	S=> E(	1197	));
			
 U1218	: Somador_Exato_1 PORT MAP(
	A=> C(	1282	),
	B=>E(	1136	),
	Cin=> Carry( 	1217	),
	Cout=> Carry( 	1218	),
	S=> E(	1198	));
			
 U1219	: Somador_Exato_1 PORT MAP(
	A=> C(	1283	),
	B=>E(	1137	),
	Cin=> Carry( 	1218	),
	Cout=> Carry( 	1219	),
	S=> E(	1199	));
			
 U1220	: Somador_Exato_1 PORT MAP(
	A=> C(	1284	),
	B=>E(	1138	),
	Cin=> Carry( 	1219	),
	Cout=> Carry( 	1220	),
	S=> E(	1200	));
			
 U1221	: Somador_Exato_1 PORT MAP(
	A=> C(	1285	),
	B=>E(	1139	),
	Cin=> Carry( 	1220	),
	Cout=> Carry( 	1221	),
	S=> E(	1201	));
			
 U1222	: Somador_Exato_1 PORT MAP(
	A=> C(	1286	),
	B=>E(	1140	),
	Cin=> Carry( 	1221	),
	Cout=> Carry( 	1222	),
	S=> E(	1202	));
			
 U1223	: Somador_Exato_1 PORT MAP(
	A=> C(	1287	),
	B=>E(	1141	),
	Cin=> Carry( 	1222	),
	Cout=> Carry( 	1223	),
	S=> E(	1203	));
			
 U1224	: Somador_Exato_1 PORT MAP(
	A=> C(	1288	),
	B=>E(	1142	),
	Cin=> Carry( 	1223	),
	Cout=> Carry( 	1224	),
	S=> E(	1204	));
			
 U1225	: Somador_Exato_1 PORT MAP(
	A=> C(	1289	),
	B=>E(	1143	),
	Cin=> Carry( 	1224	),
	Cout=> Carry( 	1225	),
	S=> E(	1205	));
			
 U1226	: Somador_Exato_1 PORT MAP(
	A=> C(	1290	),
	B=>E(	1144	),
	Cin=> Carry( 	1225	),
	Cout=> Carry( 	1226	),
	S=> E(	1206	));
			
 U1227	: Somador_Exato_1 PORT MAP(
	A=> C(	1291	),
	B=>E(	1145	),
	Cin=> Carry( 	1226	),
	Cout=> Carry( 	1227	),
	S=> E(	1207	));
			
 U1228	: Somador_Exato_1 PORT MAP(
	A=> C(	1292	),
	B=>E(	1146	),
	Cin=> Carry( 	1227	),
	Cout=> Carry( 	1228	),
	S=> E(	1208	));
			
 U1229	: Somador_Exato_1 PORT MAP(
	A=> C(	1293	),
	B=>E(	1147	),
	Cin=> Carry( 	1228	),
	Cout=> Carry( 	1229	),
	S=> E(	1209	));
			
 U1230	: Somador_Exato_1 PORT MAP(
	A=> C(	1294	),
	B=>E(	1148	),
	Cin=> Carry( 	1229	),
	Cout=> Carry( 	1230	),
	S=> E(	1210	));
			
 U1231	: Somador_Exato_1 PORT MAP(
	A=> C(	1295	),
	B=>E(	1149	),
	Cin=> Carry( 	1230	),
	Cout=> Carry( 	1231	),
	S=> E(	1211	));
			
 U1232	: Somador_Exato_1 PORT MAP(
	A=> C(	1296	),
	B=>E(	1150	),
	Cin=> Carry( 	1231	),
	Cout=> Carry( 	1232	),
	S=> E(	1212	));
			
 U1233	: Somador_Exato_1 PORT MAP(
	A=> C(	1297	),
	B=>E(	1151	),
	Cin=> Carry( 	1232	),
	Cout=> Carry( 	1233	),
	S=> E(	1213	));
			
 U1234	: Somador_Exato_1 PORT MAP(
	A=> C(	1298	),
	B=>E(	1152	),
	Cin=> Carry( 	1233	),
	Cout=> Carry( 	1234	),
	S=> E(	1214	));
			
 U1235	: Somador_Exato_1 PORT MAP(
	A=> C(	1299	),
	B=>E(	1153	),
	Cin=> Carry( 	1234	),
	Cout=> Carry( 	1235	),
	S=> E(	1215	));
			
 U1236	: Somador_Exato_1 PORT MAP(
	A=> C(	1300	),
	B=>E(	1154	),
	Cin=> Carry( 	1235	),
	Cout=> Carry( 	1236	),
	S=> E(	1216	));
			
 U1237	: Somador_Exato_1 PORT MAP(
	A=> C(	1301	),
	B=>E(	1155	),
	Cin=> Carry( 	1236	),
	Cout=> Carry( 	1237	),
	S=> E(	1217	));
			
 U1238	: Somador_Exato_1 PORT MAP(
	A=> C(	1302	),
	B=>E(	1156	),
	Cin=> Carry( 	1237	),
	Cout=> Carry( 	1238	),
	S=> E(	1218	));
			
 U1239	: Somador_Exato_1 PORT MAP(
	A=> C(	1303	),
	B=>E(	1157	),
	Cin=> Carry( 	1238	),
	Cout=> Carry( 	1239	),
	S=> E(	1219	));
			
 U1240	: Somador_Exato_1 PORT MAP(
	A=> C(	1304	),
	B=>E(	1158	),
	Cin=> Carry( 	1239	),
	Cout=> Carry( 	1240	),
	S=> E(	1220	));
			
 U1241	: Somador_Exato_1 PORT MAP(
	A=> C(	1305	),
	B=>E(	1159	),
	Cin=> Carry( 	1240	),
	Cout=> Carry( 	1241	),
	S=> E(	1221	));
			
 U1242	: Somador_Exato_1 PORT MAP(
	A=> C(	1306	),
	B=>E(	1160	),
	Cin=> Carry( 	1241	),
	Cout=> Carry( 	1242	),
	S=> E(	1222	));
			
 U1243	: Somador_Exato_1 PORT MAP(
	A=> C(	1307	),
	B=>E(	1161	),
	Cin=> Carry( 	1242	),
	Cout=> Carry( 	1243	),
	S=> E(	1223	));
			
 U1244	: Somador_Exato_1 PORT MAP(
	A=> C(	1308	),
	B=>E(	1162	),
	Cin=> Carry( 	1243	),
	Cout=> Carry( 	1244	),
	S=> E(	1224	));
			
 U1245	: Somador_Exato_1 PORT MAP(
	A=> C(	1309	),
	B=>E(	1163	),
	Cin=> Carry( 	1244	),
	Cout=> Carry( 	1245	),
	S=> E(	1225	));
			
 U1246	: Somador_Exato_1 PORT MAP(
	A=> C(	1310	),
	B=>E(	1164	),
	Cin=> Carry( 	1245	),
	Cout=> Carry( 	1246	),
	S=> E(	1226	));
			
 U1247	: Somador_Exato_1 PORT MAP(
	A=> C(	1311	),
	B=>E(	1165	),
	Cin=> Carry( 	1246	),
	Cout=> Carry( 	1247	),
	S=> E(	1227	));
			
 U1248	: Somador_Exato_1 PORT MAP(
	A=> C(	1312	),
	B=>E(	1166	),
	Cin=> Carry( 	1247	),
	Cout=> Carry( 	1248	),
	S=> E(	1228	));
			
 U1249	: Somador_Exato_1 PORT MAP(
	A=> C(	1313	),
	B=>E(	1167	),
	Cin=> Carry( 	1248	),
	Cout=> Carry( 	1249	),
	S=> E(	1229	));
			
 U1250	: Somador_Exato_1 PORT MAP(
	A=> C(	1314	),
	B=>E(	1168	),
	Cin=> Carry( 	1249	),
	Cout=> Carry( 	1250	),
	S=> E(	1230	));
			
 U1251	: Somador_Exato_1 PORT MAP(
	A=> C(	1315	),
	B=>E(	1169	),
	Cin=> Carry( 	1250	),
	Cout=> Carry( 	1251	),
	S=> E(	1231	));
			
 U1252	: Somador_Exato_1 PORT MAP(
	A=> C(	1316	),
	B=>E(	1170	),
	Cin=> Carry( 	1251	),
	Cout=> Carry( 	1252	),
	S=> E(	1232	));
			
 U1253	: Somador_Exato_1 PORT MAP(
	A=> C(	1317	),
	B=>E(	1171	),
	Cin=> Carry( 	1252	),
	Cout=> Carry( 	1253	),
	S=> E(	1233	));
			
 U1254	: Somador_Exato_1 PORT MAP(
	A=> C(	1318	),
	B=>E(	1172	),
	Cin=> Carry( 	1253	),
	Cout=> Carry( 	1254	),
	S=> E(	1234	));
			
 U1255	: Somador_Exato_1 PORT MAP(
	A=> C(	1319	),
	B=>E(	1173	),
	Cin=> Carry( 	1254	),
	Cout=> Carry( 	1255	),
	S=> E(	1235	));
			
 U1256	: Somador_Exato_1 PORT MAP(
	A=> C(	1320	),
	B=>E(	1174	),
	Cin=> Carry( 	1255	),
	Cout=> Carry( 	1256	),
	S=> E(	1236	));
			
 U1257	: Somador_Exato_1 PORT MAP(
	A=> C(	1321	),
	B=>E(	1175	),
	Cin=> Carry( 	1256	),
	Cout=> Carry( 	1257	),
	S=> E(	1237	));
			
 U1258	: Somador_Exato_1 PORT MAP(
	A=> C(	1322	),
	B=>E(	1176	),
	Cin=> Carry( 	1257	),
	Cout=> Carry( 	1258	),
	S=> E(	1238	));
			
 U1259	: Somador_Exato_1 PORT MAP(
	A=> C(	1323	),
	B=>E(	1177	),
	Cin=> Carry( 	1258	),
	Cout=> Carry( 	1259	),
	S=> E(	1239	));
			
 U1260	: Somador_Exato_1 PORT MAP(
	A=> C(	1324	),
	B=>E(	1178	),
	Cin=> Carry( 	1259	),
	Cout=> Carry( 	1260	),
	S=> E(	1240	));
			
 U1261	: Somador_Exato_1 PORT MAP(
	A=> C(	1325	),
	B=>E(	1179	),
	Cin=> Carry( 	1260	),
	Cout=> Carry( 	1261	),
	S=> E(	1241	));
			
 U1262	: Somador_Exato_1 PORT MAP(
	A=> C(	1326	),
	B=>E(	1180	),
	Cin=> Carry( 	1261	),
	Cout=> Carry( 	1262	),
	S=> E(	1242	));
			
 U1263	: Somador_Exato_1 PORT MAP(
	A=> C(	1327	),
	B=>E(	1181	),
	Cin=> Carry( 	1262	),
	Cout=> Carry( 	1263	),
	S=> E(	1243	));
			
 U1264	: Somador_Exato_1 PORT MAP(
	A=> C(	1328	),
	B=>E(	1182	),
	Cin=> Carry( 	1263	),
	Cout=> Carry( 	1264	),
	S=> E(	1244	));
			
 U1265	: Somador_Exato_1 PORT MAP(
	A=> C(	1329	),
	B=>E(	1183	),
	Cin=> Carry( 	1264	),
	Cout=> Carry( 	1265	),
	S=> E(	1245	));
			
 U1266	: Somador_Exato_1 PORT MAP(
	A=> C(	1330	),
	B=>E(	1184	),
	Cin=> Carry( 	1265	),
	Cout=> Carry( 	1266	),
	S=> E(	1246	));
			
 U1267	: Somador_Exato_1 PORT MAP(
	A=> C(	1331	),
	B=>E(	1185	),
	Cin=> Carry( 	1266	),
	Cout=> Carry( 	1267	),
	S=> E(	1247	));
			
 U1268	: Somador_Exato_1 PORT MAP(
	A=> C(	1332	),
	B=>E(	1186	),
	Cin=> Carry( 	1267	),
	Cout=> Carry( 	1268	),
	S=> E(	1248	));
			
 U1269	: Somador_Exato_1 PORT MAP(
	A=> C(	1333	),
	B=>E(	1187	),
	Cin=> Carry( 	1268	),
	Cout=> Carry( 	1269	),
	S=> E(	1249	));
			
 U1270	: Somador_Exato_1 PORT MAP(
	A=> C(	1334	),
	B=>E(	1188	),
	Cin=> Carry( 	1269	),
	Cout=> Carry( 	1270	),
	S=> E(	1250	));
			
 U1271	: Somador_Exato_1 PORT MAP(
	A=> C(	1335	),
	B=>E(	1189	),
	Cin=> Carry( 	1270	),
	Cout=> Carry( 	1271	),
	S=> E(	1251	));
			
 U1272	: Somador_Exato_1 PORT MAP(
	A=> C(	1336	),
	B=>E(	1190	),
	Cin=> Carry( 	1271	),
	Cout=> Carry( 	1272	),
	S=> E(	1252	));
			
 U1273	: Somador_Exato_1 PORT MAP(
	A=> C(	1337	),
	B=>E(	1191	),
	Cin=> Carry( 	1272	),
	Cout=> Carry( 	1273	),
	S=> E(	1253	));
			
 U1274	: Somador_Exato_1 PORT MAP(
	A=> C(	1338	),
	B=>E(	1192	),
	Cin=> Carry( 	1273	),
	Cout=> Carry( 	1274	),
	S=> E(	1254	));
			
 U1275	: Somador_Exato_1 PORT MAP(
	A=> C(	1339	),
	B=>E(	1193	),
	Cin=> Carry( 	1274	),
	Cout=> Carry( 	1275	),
	S=> E(	1255	));
			
 U1276	: Somador_Exato_1 PORT MAP(
	A=> C(	1340	),
	B=>E(	1194	),
	Cin=> Carry( 	1275	),
	Cout=> Carry( 	1276	),
	S=> E(	1256	));
			
 U1277	: Somador_Exato_1 PORT MAP(
	A=> C(	1341	),
	B=>E(	1195	),
	Cin=> Carry( 	1276	),
	Cout=> Carry( 	1277	),
	S=> E(	1257	));
			
 U1278	: Somador_Exato_1 PORT MAP(
	A=> C(	1342	),
	B=>E(	1196	),
	Cin=> Carry( 	1277	),
	Cout=> Carry( 	1278	),
	S=> E(	1258	));
			
 U1279	: Somador_Exato_1 PORT MAP(
	A=> C(	1343	),
	B=>Carry(	1215	),
	Cin=> Carry( 	1278	),
	Cout=> Carry( 	1279	),
	S=> E(	1259	));

			
 U1280	: Somador_Exato_1 PORT MAP(
	A=> C(	1344	),
	B=>E(	1197	),
	Cin=> '0'	,
	Cout=> Carry( 	1280	),
	S=> R(	21	));
			
 U1281	: Somador_Exato_1 PORT MAP(
	A=> C(	1345	),
	B=>E(	1198	),
	Cin=> Carry( 	1280	),
	Cout=> Carry( 	1281	),
	S=> E(	1260	));
			
 U1282	: Somador_Exato_1 PORT MAP(
	A=> C(	1346	),
	B=>E(	1199	),
	Cin=> Carry( 	1281	),
	Cout=> Carry( 	1282	),
	S=> E(	1261	));
			
 U1283	: Somador_Exato_1 PORT MAP(
	A=> C(	1347	),
	B=>E(	1200	),
	Cin=> Carry( 	1282	),
	Cout=> Carry( 	1283	),
	S=> E(	1262	));
			
 U1284	: Somador_Exato_1 PORT MAP(
	A=> C(	1348	),
	B=>E(	1201	),
	Cin=> Carry( 	1283	),
	Cout=> Carry( 	1284	),
	S=> E(	1263	));
			
 U1285	: Somador_Exato_1 PORT MAP(
	A=> C(	1349	),
	B=>E(	1202	),
	Cin=> Carry( 	1284	),
	Cout=> Carry( 	1285	),
	S=> E(	1264	));
			
 U1286	: Somador_Exato_1 PORT MAP(
	A=> C(	1350	),
	B=>E(	1203	),
	Cin=> Carry( 	1285	),
	Cout=> Carry( 	1286	),
	S=> E(	1265	));
			
 U1287	: Somador_Exato_1 PORT MAP(
	A=> C(	1351	),
	B=>E(	1204	),
	Cin=> Carry( 	1286	),
	Cout=> Carry( 	1287	),
	S=> E(	1266	));
			
 U1288	: Somador_Exato_1 PORT MAP(
	A=> C(	1352	),
	B=>E(	1205	),
	Cin=> Carry( 	1287	),
	Cout=> Carry( 	1288	),
	S=> E(	1267	));
			
 U1289	: Somador_Exato_1 PORT MAP(
	A=> C(	1353	),
	B=>E(	1206	),
	Cin=> Carry( 	1288	),
	Cout=> Carry( 	1289	),
	S=> E(	1268	));
			
 U1290	: Somador_Exato_1 PORT MAP(
	A=> C(	1354	),
	B=>E(	1207	),
	Cin=> Carry( 	1289	),
	Cout=> Carry( 	1290	),
	S=> E(	1269	));
			
 U1291	: Somador_Exato_1 PORT MAP(
	A=> C(	1355	),
	B=>E(	1208	),
	Cin=> Carry( 	1290	),
	Cout=> Carry( 	1291	),
	S=> E(	1270	));
			
 U1292	: Somador_Exato_1 PORT MAP(
	A=> C(	1356	),
	B=>E(	1209	),
	Cin=> Carry( 	1291	),
	Cout=> Carry( 	1292	),
	S=> E(	1271	));
			
 U1293	: Somador_Exato_1 PORT MAP(
	A=> C(	1357	),
	B=>E(	1210	),
	Cin=> Carry( 	1292	),
	Cout=> Carry( 	1293	),
	S=> E(	1272	));
			
 U1294	: Somador_Exato_1 PORT MAP(
	A=> C(	1358	),
	B=>E(	1211	),
	Cin=> Carry( 	1293	),
	Cout=> Carry( 	1294	),
	S=> E(	1273	));
			
 U1295	: Somador_Exato_1 PORT MAP(
	A=> C(	1359	),
	B=>E(	1212	),
	Cin=> Carry( 	1294	),
	Cout=> Carry( 	1295	),
	S=> E(	1274	));
			
 U1296	: Somador_Exato_1 PORT MAP(
	A=> C(	1360	),
	B=>E(	1213	),
	Cin=> Carry( 	1295	),
	Cout=> Carry( 	1296	),
	S=> E(	1275	));
			
 U1297	: Somador_Exato_1 PORT MAP(
	A=> C(	1361	),
	B=>E(	1214	),
	Cin=> Carry( 	1296	),
	Cout=> Carry( 	1297	),
	S=> E(	1276	));
			
 U1298	: Somador_Exato_1 PORT MAP(
	A=> C(	1362	),
	B=>E(	1215	),
	Cin=> Carry( 	1297	),
	Cout=> Carry( 	1298	),
	S=> E(	1277	));
			
 U1299	: Somador_Exato_1 PORT MAP(
	A=> C(	1363	),
	B=>E(	1216	),
	Cin=> Carry( 	1298	),
	Cout=> Carry( 	1299	),
	S=> E(	1278	));
			
 U1300	: Somador_Exato_1 PORT MAP(
	A=> C(	1364	),
	B=>E(	1217	),
	Cin=> Carry( 	1299	),
	Cout=> Carry( 	1300	),
	S=> E(	1279	));
			
 U1301	: Somador_Exato_1 PORT MAP(
	A=> C(	1365	),
	B=>E(	1218	),
	Cin=> Carry( 	1300	),
	Cout=> Carry( 	1301	),
	S=> E(	1280	));
			
 U1302	: Somador_Exato_1 PORT MAP(
	A=> C(	1366	),
	B=>E(	1219	),
	Cin=> Carry( 	1301	),
	Cout=> Carry( 	1302	),
	S=> E(	1281	));
			
 U1303	: Somador_Exato_1 PORT MAP(
	A=> C(	1367	),
	B=>E(	1220	),
	Cin=> Carry( 	1302	),
	Cout=> Carry( 	1303	),
	S=> E(	1282	));
			
 U1304	: Somador_Exato_1 PORT MAP(
	A=> C(	1368	),
	B=>E(	1221	),
	Cin=> Carry( 	1303	),
	Cout=> Carry( 	1304	),
	S=> E(	1283	));
			
 U1305	: Somador_Exato_1 PORT MAP(
	A=> C(	1369	),
	B=>E(	1222	),
	Cin=> Carry( 	1304	),
	Cout=> Carry( 	1305	),
	S=> E(	1284	));
			
 U1306	: Somador_Exato_1 PORT MAP(
	A=> C(	1370	),
	B=>E(	1223	),
	Cin=> Carry( 	1305	),
	Cout=> Carry( 	1306	),
	S=> E(	1285	));
			
 U1307	: Somador_Exato_1 PORT MAP(
	A=> C(	1371	),
	B=>E(	1224	),
	Cin=> Carry( 	1306	),
	Cout=> Carry( 	1307	),
	S=> E(	1286	));
			
 U1308	: Somador_Exato_1 PORT MAP(
	A=> C(	1372	),
	B=>E(	1225	),
	Cin=> Carry( 	1307	),
	Cout=> Carry( 	1308	),
	S=> E(	1287	));
			
 U1309	: Somador_Exato_1 PORT MAP(
	A=> C(	1373	),
	B=>E(	1226	),
	Cin=> Carry( 	1308	),
	Cout=> Carry( 	1309	),
	S=> E(	1288	));
			
 U1310	: Somador_Exato_1 PORT MAP(
	A=> C(	1374	),
	B=>E(	1227	),
	Cin=> Carry( 	1309	),
	Cout=> Carry( 	1310	),
	S=> E(	1289	));
			
 U1311	: Somador_Exato_1 PORT MAP(
	A=> C(	1375	),
	B=>E(	1228	),
	Cin=> Carry( 	1310	),
	Cout=> Carry( 	1311	),
	S=> E(	1290	));
			
 U1312	: Somador_Exato_1 PORT MAP(
	A=> C(	1376	),
	B=>E(	1229	),
	Cin=> Carry( 	1311	),
	Cout=> Carry( 	1312	),
	S=> E(	1291	));
			
 U1313	: Somador_Exato_1 PORT MAP(
	A=> C(	1377	),
	B=>E(	1230	),
	Cin=> Carry( 	1312	),
	Cout=> Carry( 	1313	),
	S=> E(	1292	));
			
 U1314	: Somador_Exato_1 PORT MAP(
	A=> C(	1378	),
	B=>E(	1231	),
	Cin=> Carry( 	1313	),
	Cout=> Carry( 	1314	),
	S=> E(	1293	));
			
 U1315	: Somador_Exato_1 PORT MAP(
	A=> C(	1379	),
	B=>E(	1232	),
	Cin=> Carry( 	1314	),
	Cout=> Carry( 	1315	),
	S=> E(	1294	));
			
 U1316	: Somador_Exato_1 PORT MAP(
	A=> C(	1380	),
	B=>E(	1233	),
	Cin=> Carry( 	1315	),
	Cout=> Carry( 	1316	),
	S=> E(	1295	));
			
 U1317	: Somador_Exato_1 PORT MAP(
	A=> C(	1381	),
	B=>E(	1234	),
	Cin=> Carry( 	1316	),
	Cout=> Carry( 	1317	),
	S=> E(	1296	));
			
 U1318	: Somador_Exato_1 PORT MAP(
	A=> C(	1382	),
	B=>E(	1235	),
	Cin=> Carry( 	1317	),
	Cout=> Carry( 	1318	),
	S=> E(	1297	));
			
 U1319	: Somador_Exato_1 PORT MAP(
	A=> C(	1383	),
	B=>E(	1236	),
	Cin=> Carry( 	1318	),
	Cout=> Carry( 	1319	),
	S=> E(	1298	));
			
 U1320	: Somador_Exato_1 PORT MAP(
	A=> C(	1384	),
	B=>E(	1237	),
	Cin=> Carry( 	1319	),
	Cout=> Carry( 	1320	),
	S=> E(	1299	));
			
 U1321	: Somador_Exato_1 PORT MAP(
	A=> C(	1385	),
	B=>E(	1238	),
	Cin=> Carry( 	1320	),
	Cout=> Carry( 	1321	),
	S=> E(	1300	));
			
 U1322	: Somador_Exato_1 PORT MAP(
	A=> C(	1386	),
	B=>E(	1239	),
	Cin=> Carry( 	1321	),
	Cout=> Carry( 	1322	),
	S=> E(	1301	));
			
 U1323	: Somador_Exato_1 PORT MAP(
	A=> C(	1387	),
	B=>E(	1240	),
	Cin=> Carry( 	1322	),
	Cout=> Carry( 	1323	),
	S=> E(	1302	));
			
 U1324	: Somador_Exato_1 PORT MAP(
	A=> C(	1388	),
	B=>E(	1241	),
	Cin=> Carry( 	1323	),
	Cout=> Carry( 	1324	),
	S=> E(	1303	));
			
 U1325	: Somador_Exato_1 PORT MAP(
	A=> C(	1389	),
	B=>E(	1242	),
	Cin=> Carry( 	1324	),
	Cout=> Carry( 	1325	),
	S=> E(	1304	));
			
 U1326	: Somador_Exato_1 PORT MAP(
	A=> C(	1390	),
	B=>E(	1243	),
	Cin=> Carry( 	1325	),
	Cout=> Carry( 	1326	),
	S=> E(	1305	));
			
 U1327	: Somador_Exato_1 PORT MAP(
	A=> C(	1391	),
	B=>E(	1244	),
	Cin=> Carry( 	1326	),
	Cout=> Carry( 	1327	),
	S=> E(	1306	));
			
 U1328	: Somador_Exato_1 PORT MAP(
	A=> C(	1392	),
	B=>E(	1245	),
	Cin=> Carry( 	1327	),
	Cout=> Carry( 	1328	),
	S=> E(	1307	));
			
 U1329	: Somador_Exato_1 PORT MAP(
	A=> C(	1393	),
	B=>E(	1246	),
	Cin=> Carry( 	1328	),
	Cout=> Carry( 	1329	),
	S=> E(	1308	));
			
 U1330	: Somador_Exato_1 PORT MAP(
	A=> C(	1394	),
	B=>E(	1247	),
	Cin=> Carry( 	1329	),
	Cout=> Carry( 	1330	),
	S=> E(	1309	));
			
 U1331	: Somador_Exato_1 PORT MAP(
	A=> C(	1395	),
	B=>E(	1248	),
	Cin=> Carry( 	1330	),
	Cout=> Carry( 	1331	),
	S=> E(	1310	));
			
 U1332	: Somador_Exato_1 PORT MAP(
	A=> C(	1396	),
	B=>E(	1249	),
	Cin=> Carry( 	1331	),
	Cout=> Carry( 	1332	),
	S=> E(	1311	));
			
 U1333	: Somador_Exato_1 PORT MAP(
	A=> C(	1397	),
	B=>E(	1250	),
	Cin=> Carry( 	1332	),
	Cout=> Carry( 	1333	),
	S=> E(	1312	));
			
 U1334	: Somador_Exato_1 PORT MAP(
	A=> C(	1398	),
	B=>E(	1251	),
	Cin=> Carry( 	1333	),
	Cout=> Carry( 	1334	),
	S=> E(	1313	));
			
 U1335	: Somador_Exato_1 PORT MAP(
	A=> C(	1399	),
	B=>E(	1252	),
	Cin=> Carry( 	1334	),
	Cout=> Carry( 	1335	),
	S=> E(	1314	));
			
 U1336	: Somador_Exato_1 PORT MAP(
	A=> C(	1400	),
	B=>E(	1253	),
	Cin=> Carry( 	1335	),
	Cout=> Carry( 	1336	),
	S=> E(	1315	));
			
 U1337	: Somador_Exato_1 PORT MAP(
	A=> C(	1401	),
	B=>E(	1254	),
	Cin=> Carry( 	1336	),
	Cout=> Carry( 	1337	),
	S=> E(	1316	));
			
 U1338	: Somador_Exato_1 PORT MAP(
	A=> C(	1402	),
	B=>E(	1255	),
	Cin=> Carry( 	1337	),
	Cout=> Carry( 	1338	),
	S=> E(	1317	));
			
 U1339	: Somador_Exato_1 PORT MAP(
	A=> C(	1403	),
	B=>E(	1256	),
	Cin=> Carry( 	1338	),
	Cout=> Carry( 	1339	),
	S=> E(	1318	));
			
 U1340	: Somador_Exato_1 PORT MAP(
	A=> C(	1404	),
	B=>E(	1257	),
	Cin=> Carry( 	1339	),
	Cout=> Carry( 	1340	),
	S=> E(	1319	));
			
 U1341	: Somador_Exato_1 PORT MAP(
	A=> C(	1405	),
	B=>E(	1258	),
	Cin=> Carry( 	1340	),
	Cout=> Carry( 	1341	),
	S=> E(	1320	));
			
 U1342	: Somador_Exato_1 PORT MAP(
	A=> C(	1406	),
	B=>E(	1259	),
	Cin=> Carry( 	1341	),
	Cout=> Carry( 	1342	),
	S=> E(	1321	));
			
 U1343	: Somador_Exato_1 PORT MAP(
	A=> C(	1407	),
	B=>Carry(	1279	),
	Cin=> Carry( 	1342	),
	Cout=> Carry( 	1343	),
	S=> E(	1322	));

			
 U1344	: Somador_Exato_1 PORT MAP(
	A=> C(	1408	),
	B=>E(	1260	),
	Cin=> '0'	,
	Cout=> Carry( 	1344	),
	S=> R(	22	));
			
 U1345	: Somador_Exato_1 PORT MAP(
	A=> C(	1409	),
	B=>E(	1261	),
	Cin=> Carry( 	1344	),
	Cout=> Carry( 	1345	),
	S=> E(	1323	));
			
 U1346	: Somador_Exato_1 PORT MAP(
	A=> C(	1410	),
	B=>E(	1262	),
	Cin=> Carry( 	1345	),
	Cout=> Carry( 	1346	),
	S=> E(	1324	));
			
 U1347	: Somador_Exato_1 PORT MAP(
	A=> C(	1411	),
	B=>E(	1263	),
	Cin=> Carry( 	1346	),
	Cout=> Carry( 	1347	),
	S=> E(	1325	));
			
 U1348	: Somador_Exato_1 PORT MAP(
	A=> C(	1412	),
	B=>E(	1264	),
	Cin=> Carry( 	1347	),
	Cout=> Carry( 	1348	),
	S=> E(	1326	));
			
 U1349	: Somador_Exato_1 PORT MAP(
	A=> C(	1413	),
	B=>E(	1265	),
	Cin=> Carry( 	1348	),
	Cout=> Carry( 	1349	),
	S=> E(	1327	));
			
 U1350	: Somador_Exato_1 PORT MAP(
	A=> C(	1414	),
	B=>E(	1266	),
	Cin=> Carry( 	1349	),
	Cout=> Carry( 	1350	),
	S=> E(	1328	));
			
 U1351	: Somador_Exato_1 PORT MAP(
	A=> C(	1415	),
	B=>E(	1267	),
	Cin=> Carry( 	1350	),
	Cout=> Carry( 	1351	),
	S=> E(	1329	));
			
 U1352	: Somador_Exato_1 PORT MAP(
	A=> C(	1416	),
	B=>E(	1268	),
	Cin=> Carry( 	1351	),
	Cout=> Carry( 	1352	),
	S=> E(	1330	));
			
 U1353	: Somador_Exato_1 PORT MAP(
	A=> C(	1417	),
	B=>E(	1269	),
	Cin=> Carry( 	1352	),
	Cout=> Carry( 	1353	),
	S=> E(	1331	));
			
 U1354	: Somador_Exato_1 PORT MAP(
	A=> C(	1418	),
	B=>E(	1270	),
	Cin=> Carry( 	1353	),
	Cout=> Carry( 	1354	),
	S=> E(	1332	));
			
 U1355	: Somador_Exato_1 PORT MAP(
	A=> C(	1419	),
	B=>E(	1271	),
	Cin=> Carry( 	1354	),
	Cout=> Carry( 	1355	),
	S=> E(	1333	));
			
 U1356	: Somador_Exato_1 PORT MAP(
	A=> C(	1420	),
	B=>E(	1272	),
	Cin=> Carry( 	1355	),
	Cout=> Carry( 	1356	),
	S=> E(	1334	));
			
 U1357	: Somador_Exato_1 PORT MAP(
	A=> C(	1421	),
	B=>E(	1273	),
	Cin=> Carry( 	1356	),
	Cout=> Carry( 	1357	),
	S=> E(	1335	));
			
 U1358	: Somador_Exato_1 PORT MAP(
	A=> C(	1422	),
	B=>E(	1274	),
	Cin=> Carry( 	1357	),
	Cout=> Carry( 	1358	),
	S=> E(	1336	));
			
 U1359	: Somador_Exato_1 PORT MAP(
	A=> C(	1423	),
	B=>E(	1275	),
	Cin=> Carry( 	1358	),
	Cout=> Carry( 	1359	),
	S=> E(	1337	));
			
 U1360	: Somador_Exato_1 PORT MAP(
	A=> C(	1424	),
	B=>E(	1276	),
	Cin=> Carry( 	1359	),
	Cout=> Carry( 	1360	),
	S=> E(	1338	));
			
 U1361	: Somador_Exato_1 PORT MAP(
	A=> C(	1425	),
	B=>E(	1277	),
	Cin=> Carry( 	1360	),
	Cout=> Carry( 	1361	),
	S=> E(	1339	));
			
 U1362	: Somador_Exato_1 PORT MAP(
	A=> C(	1426	),
	B=>E(	1278	),
	Cin=> Carry( 	1361	),
	Cout=> Carry( 	1362	),
	S=> E(	1340	));
			
 U1363	: Somador_Exato_1 PORT MAP(
	A=> C(	1427	),
	B=>E(	1279	),
	Cin=> Carry( 	1362	),
	Cout=> Carry( 	1363	),
	S=> E(	1341	));
			
 U1364	: Somador_Exato_1 PORT MAP(
	A=> C(	1428	),
	B=>E(	1280	),
	Cin=> Carry( 	1363	),
	Cout=> Carry( 	1364	),
	S=> E(	1342	));
			
 U1365	: Somador_Exato_1 PORT MAP(
	A=> C(	1429	),
	B=>E(	1281	),
	Cin=> Carry( 	1364	),
	Cout=> Carry( 	1365	),
	S=> E(	1343	));
			
 U1366	: Somador_Exato_1 PORT MAP(
	A=> C(	1430	),
	B=>E(	1282	),
	Cin=> Carry( 	1365	),
	Cout=> Carry( 	1366	),
	S=> E(	1344	));
			
 U1367	: Somador_Exato_1 PORT MAP(
	A=> C(	1431	),
	B=>E(	1283	),
	Cin=> Carry( 	1366	),
	Cout=> Carry( 	1367	),
	S=> E(	1345	));
			
 U1368	: Somador_Exato_1 PORT MAP(
	A=> C(	1432	),
	B=>E(	1284	),
	Cin=> Carry( 	1367	),
	Cout=> Carry( 	1368	),
	S=> E(	1346	));
			
 U1369	: Somador_Exato_1 PORT MAP(
	A=> C(	1433	),
	B=>E(	1285	),
	Cin=> Carry( 	1368	),
	Cout=> Carry( 	1369	),
	S=> E(	1347	));
			
 U1370	: Somador_Exato_1 PORT MAP(
	A=> C(	1434	),
	B=>E(	1286	),
	Cin=> Carry( 	1369	),
	Cout=> Carry( 	1370	),
	S=> E(	1348	));
			
 U1371	: Somador_Exato_1 PORT MAP(
	A=> C(	1435	),
	B=>E(	1287	),
	Cin=> Carry( 	1370	),
	Cout=> Carry( 	1371	),
	S=> E(	1349	));
			
 U1372	: Somador_Exato_1 PORT MAP(
	A=> C(	1436	),
	B=>E(	1288	),
	Cin=> Carry( 	1371	),
	Cout=> Carry( 	1372	),
	S=> E(	1350	));
			
 U1373	: Somador_Exato_1 PORT MAP(
	A=> C(	1437	),
	B=>E(	1289	),
	Cin=> Carry( 	1372	),
	Cout=> Carry( 	1373	),
	S=> E(	1351	));
			
 U1374	: Somador_Exato_1 PORT MAP(
	A=> C(	1438	),
	B=>E(	1290	),
	Cin=> Carry( 	1373	),
	Cout=> Carry( 	1374	),
	S=> E(	1352	));
			
 U1375	: Somador_Exato_1 PORT MAP(
	A=> C(	1439	),
	B=>E(	1291	),
	Cin=> Carry( 	1374	),
	Cout=> Carry( 	1375	),
	S=> E(	1353	));
			
 U1376	: Somador_Exato_1 PORT MAP(
	A=> C(	1440	),
	B=>E(	1292	),
	Cin=> Carry( 	1375	),
	Cout=> Carry( 	1376	),
	S=> E(	1354	));
			
 U1377	: Somador_Exato_1 PORT MAP(
	A=> C(	1441	),
	B=>E(	1293	),
	Cin=> Carry( 	1376	),
	Cout=> Carry( 	1377	),
	S=> E(	1355	));
			
 U1378	: Somador_Exato_1 PORT MAP(
	A=> C(	1442	),
	B=>E(	1294	),
	Cin=> Carry( 	1377	),
	Cout=> Carry( 	1378	),
	S=> E(	1356	));
			
 U1379	: Somador_Exato_1 PORT MAP(
	A=> C(	1443	),
	B=>E(	1295	),
	Cin=> Carry( 	1378	),
	Cout=> Carry( 	1379	),
	S=> E(	1357	));
			
 U1380	: Somador_Exato_1 PORT MAP(
	A=> C(	1444	),
	B=>E(	1296	),
	Cin=> Carry( 	1379	),
	Cout=> Carry( 	1380	),
	S=> E(	1358	));
			
 U1381	: Somador_Exato_1 PORT MAP(
	A=> C(	1445	),
	B=>E(	1297	),
	Cin=> Carry( 	1380	),
	Cout=> Carry( 	1381	),
	S=> E(	1359	));
			
 U1382	: Somador_Exato_1 PORT MAP(
	A=> C(	1446	),
	B=>E(	1298	),
	Cin=> Carry( 	1381	),
	Cout=> Carry( 	1382	),
	S=> E(	1360	));
			
 U1383	: Somador_Exato_1 PORT MAP(
	A=> C(	1447	),
	B=>E(	1299	),
	Cin=> Carry( 	1382	),
	Cout=> Carry( 	1383	),
	S=> E(	1361	));
			
 U1384	: Somador_Exato_1 PORT MAP(
	A=> C(	1448	),
	B=>E(	1300	),
	Cin=> Carry( 	1383	),
	Cout=> Carry( 	1384	),
	S=> E(	1362	));
			
 U1385	: Somador_Exato_1 PORT MAP(
	A=> C(	1449	),
	B=>E(	1301	),
	Cin=> Carry( 	1384	),
	Cout=> Carry( 	1385	),
	S=> E(	1363	));
			
 U1386	: Somador_Exato_1 PORT MAP(
	A=> C(	1450	),
	B=>E(	1302	),
	Cin=> Carry( 	1385	),
	Cout=> Carry( 	1386	),
	S=> E(	1364	));
			
 U1387	: Somador_Exato_1 PORT MAP(
	A=> C(	1451	),
	B=>E(	1303	),
	Cin=> Carry( 	1386	),
	Cout=> Carry( 	1387	),
	S=> E(	1365	));
			
 U1388	: Somador_Exato_1 PORT MAP(
	A=> C(	1452	),
	B=>E(	1304	),
	Cin=> Carry( 	1387	),
	Cout=> Carry( 	1388	),
	S=> E(	1366	));
			
 U1389	: Somador_Exato_1 PORT MAP(
	A=> C(	1453	),
	B=>E(	1305	),
	Cin=> Carry( 	1388	),
	Cout=> Carry( 	1389	),
	S=> E(	1367	));
			
 U1390	: Somador_Exato_1 PORT MAP(
	A=> C(	1454	),
	B=>E(	1306	),
	Cin=> Carry( 	1389	),
	Cout=> Carry( 	1390	),
	S=> E(	1368	));
			
 U1391	: Somador_Exato_1 PORT MAP(
	A=> C(	1455	),
	B=>E(	1307	),
	Cin=> Carry( 	1390	),
	Cout=> Carry( 	1391	),
	S=> E(	1369	));
			
 U1392	: Somador_Exato_1 PORT MAP(
	A=> C(	1456	),
	B=>E(	1308	),
	Cin=> Carry( 	1391	),
	Cout=> Carry( 	1392	),
	S=> E(	1370	));
			
 U1393	: Somador_Exato_1 PORT MAP(
	A=> C(	1457	),
	B=>E(	1309	),
	Cin=> Carry( 	1392	),
	Cout=> Carry( 	1393	),
	S=> E(	1371	));
			
 U1394	: Somador_Exato_1 PORT MAP(
	A=> C(	1458	),
	B=>E(	1310	),
	Cin=> Carry( 	1393	),
	Cout=> Carry( 	1394	),
	S=> E(	1372	));
			
 U1395	: Somador_Exato_1 PORT MAP(
	A=> C(	1459	),
	B=>E(	1311	),
	Cin=> Carry( 	1394	),
	Cout=> Carry( 	1395	),
	S=> E(	1373	));
			
 U1396	: Somador_Exato_1 PORT MAP(
	A=> C(	1460	),
	B=>E(	1312	),
	Cin=> Carry( 	1395	),
	Cout=> Carry( 	1396	),
	S=> E(	1374	));
			
 U1397	: Somador_Exato_1 PORT MAP(
	A=> C(	1461	),
	B=>E(	1313	),
	Cin=> Carry( 	1396	),
	Cout=> Carry( 	1397	),
	S=> E(	1375	));
			
 U1398	: Somador_Exato_1 PORT MAP(
	A=> C(	1462	),
	B=>E(	1314	),
	Cin=> Carry( 	1397	),
	Cout=> Carry( 	1398	),
	S=> E(	1376	));
			
 U1399	: Somador_Exato_1 PORT MAP(
	A=> C(	1463	),
	B=>E(	1315	),
	Cin=> Carry( 	1398	),
	Cout=> Carry( 	1399	),
	S=> E(	1377	));
			
 U1400	: Somador_Exato_1 PORT MAP(
	A=> C(	1464	),
	B=>E(	1316	),
	Cin=> Carry( 	1399	),
	Cout=> Carry( 	1400	),
	S=> E(	1378	));
			
 U1401	: Somador_Exato_1 PORT MAP(
	A=> C(	1465	),
	B=>E(	1317	),
	Cin=> Carry( 	1400	),
	Cout=> Carry( 	1401	),
	S=> E(	1379	));
			
 U1402	: Somador_Exato_1 PORT MAP(
	A=> C(	1466	),
	B=>E(	1318	),
	Cin=> Carry( 	1401	),
	Cout=> Carry( 	1402	),
	S=> E(	1380	));
			
 U1403	: Somador_Exato_1 PORT MAP(
	A=> C(	1467	),
	B=>E(	1319	),
	Cin=> Carry( 	1402	),
	Cout=> Carry( 	1403	),
	S=> E(	1381	));
			
 U1404	: Somador_Exato_1 PORT MAP(
	A=> C(	1468	),
	B=>E(	1320	),
	Cin=> Carry( 	1403	),
	Cout=> Carry( 	1404	),
	S=> E(	1382	));
			
 U1405	: Somador_Exato_1 PORT MAP(
	A=> C(	1469	),
	B=>E(	1321	),
	Cin=> Carry( 	1404	),
	Cout=> Carry( 	1405	),
	S=> E(	1383	));
			
 U1406	: Somador_Exato_1 PORT MAP(
	A=> C(	1470	),
	B=>E(	1322	),
	Cin=> Carry( 	1405	),
	Cout=> Carry( 	1406	),
	S=> E(	1384	));
			
 U1407	: Somador_Exato_1 PORT MAP(
	A=> C(	1471	),
	B=>Carry(	1343	),
	Cin=> Carry( 	1406	),
	Cout=> Carry( 	1407	),
	S=> E(	1385	));

			
 U1408	: Somador_Exato_1 PORT MAP(
	A=> C(	1472	),
	B=>E(	1323	),
	Cin=> '0'	,
	Cout=> Carry( 	1408	),
	S=> R(	23	));
			
 U1409	: Somador_Exato_1 PORT MAP(
	A=> C(	1473	),
	B=>E(	1324	),
	Cin=> Carry( 	1408	),
	Cout=> Carry( 	1409	),
	S=> E(	1386	));
			
 U1410	: Somador_Exato_1 PORT MAP(
	A=> C(	1474	),
	B=>E(	1325	),
	Cin=> Carry( 	1409	),
	Cout=> Carry( 	1410	),
	S=> E(	1387	));
			
 U1411	: Somador_Exato_1 PORT MAP(
	A=> C(	1475	),
	B=>E(	1326	),
	Cin=> Carry( 	1410	),
	Cout=> Carry( 	1411	),
	S=> E(	1388	));
			
 U1412	: Somador_Exato_1 PORT MAP(
	A=> C(	1476	),
	B=>E(	1327	),
	Cin=> Carry( 	1411	),
	Cout=> Carry( 	1412	),
	S=> E(	1389	));
			
 U1413	: Somador_Exato_1 PORT MAP(
	A=> C(	1477	),
	B=>E(	1328	),
	Cin=> Carry( 	1412	),
	Cout=> Carry( 	1413	),
	S=> E(	1390	));
			
 U1414	: Somador_Exato_1 PORT MAP(
	A=> C(	1478	),
	B=>E(	1329	),
	Cin=> Carry( 	1413	),
	Cout=> Carry( 	1414	),
	S=> E(	1391	));
			
 U1415	: Somador_Exato_1 PORT MAP(
	A=> C(	1479	),
	B=>E(	1330	),
	Cin=> Carry( 	1414	),
	Cout=> Carry( 	1415	),
	S=> E(	1392	));
			
 U1416	: Somador_Exato_1 PORT MAP(
	A=> C(	1480	),
	B=>E(	1331	),
	Cin=> Carry( 	1415	),
	Cout=> Carry( 	1416	),
	S=> E(	1393	));
			
 U1417	: Somador_Exato_1 PORT MAP(
	A=> C(	1481	),
	B=>E(	1332	),
	Cin=> Carry( 	1416	),
	Cout=> Carry( 	1417	),
	S=> E(	1394	));
			
 U1418	: Somador_Exato_1 PORT MAP(
	A=> C(	1482	),
	B=>E(	1333	),
	Cin=> Carry( 	1417	),
	Cout=> Carry( 	1418	),
	S=> E(	1395	));
			
 U1419	: Somador_Exato_1 PORT MAP(
	A=> C(	1483	),
	B=>E(	1334	),
	Cin=> Carry( 	1418	),
	Cout=> Carry( 	1419	),
	S=> E(	1396	));
			
 U1420	: Somador_Exato_1 PORT MAP(
	A=> C(	1484	),
	B=>E(	1335	),
	Cin=> Carry( 	1419	),
	Cout=> Carry( 	1420	),
	S=> E(	1397	));
			
 U1421	: Somador_Exato_1 PORT MAP(
	A=> C(	1485	),
	B=>E(	1336	),
	Cin=> Carry( 	1420	),
	Cout=> Carry( 	1421	),
	S=> E(	1398	));
			
 U1422	: Somador_Exato_1 PORT MAP(
	A=> C(	1486	),
	B=>E(	1337	),
	Cin=> Carry( 	1421	),
	Cout=> Carry( 	1422	),
	S=> E(	1399	));
			
 U1423	: Somador_Exato_1 PORT MAP(
	A=> C(	1487	),
	B=>E(	1338	),
	Cin=> Carry( 	1422	),
	Cout=> Carry( 	1423	),
	S=> E(	1400	));
			
 U1424	: Somador_Exato_1 PORT MAP(
	A=> C(	1488	),
	B=>E(	1339	),
	Cin=> Carry( 	1423	),
	Cout=> Carry( 	1424	),
	S=> E(	1401	));
			
 U1425	: Somador_Exato_1 PORT MAP(
	A=> C(	1489	),
	B=>E(	1340	),
	Cin=> Carry( 	1424	),
	Cout=> Carry( 	1425	),
	S=> E(	1402	));
			
 U1426	: Somador_Exato_1 PORT MAP(
	A=> C(	1490	),
	B=>E(	1341	),
	Cin=> Carry( 	1425	),
	Cout=> Carry( 	1426	),
	S=> E(	1403	));
			
 U1427	: Somador_Exato_1 PORT MAP(
	A=> C(	1491	),
	B=>E(	1342	),
	Cin=> Carry( 	1426	),
	Cout=> Carry( 	1427	),
	S=> E(	1404	));
			
 U1428	: Somador_Exato_1 PORT MAP(
	A=> C(	1492	),
	B=>E(	1343	),
	Cin=> Carry( 	1427	),
	Cout=> Carry( 	1428	),
	S=> E(	1405	));
			
 U1429	: Somador_Exato_1 PORT MAP(
	A=> C(	1493	),
	B=>E(	1344	),
	Cin=> Carry( 	1428	),
	Cout=> Carry( 	1429	),
	S=> E(	1406	));
			
 U1430	: Somador_Exato_1 PORT MAP(
	A=> C(	1494	),
	B=>E(	1345	),
	Cin=> Carry( 	1429	),
	Cout=> Carry( 	1430	),
	S=> E(	1407	));
			
 U1431	: Somador_Exato_1 PORT MAP(
	A=> C(	1495	),
	B=>E(	1346	),
	Cin=> Carry( 	1430	),
	Cout=> Carry( 	1431	),
	S=> E(	1408	));
			
 U1432	: Somador_Exato_1 PORT MAP(
	A=> C(	1496	),
	B=>E(	1347	),
	Cin=> Carry( 	1431	),
	Cout=> Carry( 	1432	),
	S=> E(	1409	));
			
 U1433	: Somador_Exato_1 PORT MAP(
	A=> C(	1497	),
	B=>E(	1348	),
	Cin=> Carry( 	1432	),
	Cout=> Carry( 	1433	),
	S=> E(	1410	));
			
 U1434	: Somador_Exato_1 PORT MAP(
	A=> C(	1498	),
	B=>E(	1349	),
	Cin=> Carry( 	1433	),
	Cout=> Carry( 	1434	),
	S=> E(	1411	));
			
 U1435	: Somador_Exato_1 PORT MAP(
	A=> C(	1499	),
	B=>E(	1350	),
	Cin=> Carry( 	1434	),
	Cout=> Carry( 	1435	),
	S=> E(	1412	));
			
 U1436	: Somador_Exato_1 PORT MAP(
	A=> C(	1500	),
	B=>E(	1351	),
	Cin=> Carry( 	1435	),
	Cout=> Carry( 	1436	),
	S=> E(	1413	));
			
 U1437	: Somador_Exato_1 PORT MAP(
	A=> C(	1501	),
	B=>E(	1352	),
	Cin=> Carry( 	1436	),
	Cout=> Carry( 	1437	),
	S=> E(	1414	));
			
 U1438	: Somador_Exato_1 PORT MAP(
	A=> C(	1502	),
	B=>E(	1353	),
	Cin=> Carry( 	1437	),
	Cout=> Carry( 	1438	),
	S=> E(	1415	));
			
 U1439	: Somador_Exato_1 PORT MAP(
	A=> C(	1503	),
	B=>E(	1354	),
	Cin=> Carry( 	1438	),
	Cout=> Carry( 	1439	),
	S=> E(	1416	));
			
 U1440	: Somador_Exato_1 PORT MAP(
	A=> C(	1504	),
	B=>E(	1355	),
	Cin=> Carry( 	1439	),
	Cout=> Carry( 	1440	),
	S=> E(	1417	));
			
 U1441	: Somador_Exato_1 PORT MAP(
	A=> C(	1505	),
	B=>E(	1356	),
	Cin=> Carry( 	1440	),
	Cout=> Carry( 	1441	),
	S=> E(	1418	));
			
 U1442	: Somador_Exato_1 PORT MAP(
	A=> C(	1506	),
	B=>E(	1357	),
	Cin=> Carry( 	1441	),
	Cout=> Carry( 	1442	),
	S=> E(	1419	));
			
 U1443	: Somador_Exato_1 PORT MAP(
	A=> C(	1507	),
	B=>E(	1358	),
	Cin=> Carry( 	1442	),
	Cout=> Carry( 	1443	),
	S=> E(	1420	));
			
 U1444	: Somador_Exato_1 PORT MAP(
	A=> C(	1508	),
	B=>E(	1359	),
	Cin=> Carry( 	1443	),
	Cout=> Carry( 	1444	),
	S=> E(	1421	));
			
 U1445	: Somador_Exato_1 PORT MAP(
	A=> C(	1509	),
	B=>E(	1360	),
	Cin=> Carry( 	1444	),
	Cout=> Carry( 	1445	),
	S=> E(	1422	));
			
 U1446	: Somador_Exato_1 PORT MAP(
	A=> C(	1510	),
	B=>E(	1361	),
	Cin=> Carry( 	1445	),
	Cout=> Carry( 	1446	),
	S=> E(	1423	));
			
 U1447	: Somador_Exato_1 PORT MAP(
	A=> C(	1511	),
	B=>E(	1362	),
	Cin=> Carry( 	1446	),
	Cout=> Carry( 	1447	),
	S=> E(	1424	));
			
 U1448	: Somador_Exato_1 PORT MAP(
	A=> C(	1512	),
	B=>E(	1363	),
	Cin=> Carry( 	1447	),
	Cout=> Carry( 	1448	),
	S=> E(	1425	));
			
 U1449	: Somador_Exato_1 PORT MAP(
	A=> C(	1513	),
	B=>E(	1364	),
	Cin=> Carry( 	1448	),
	Cout=> Carry( 	1449	),
	S=> E(	1426	));
			
 U1450	: Somador_Exato_1 PORT MAP(
	A=> C(	1514	),
	B=>E(	1365	),
	Cin=> Carry( 	1449	),
	Cout=> Carry( 	1450	),
	S=> E(	1427	));
			
 U1451	: Somador_Exato_1 PORT MAP(
	A=> C(	1515	),
	B=>E(	1366	),
	Cin=> Carry( 	1450	),
	Cout=> Carry( 	1451	),
	S=> E(	1428	));
			
 U1452	: Somador_Exato_1 PORT MAP(
	A=> C(	1516	),
	B=>E(	1367	),
	Cin=> Carry( 	1451	),
	Cout=> Carry( 	1452	),
	S=> E(	1429	));
			
 U1453	: Somador_Exato_1 PORT MAP(
	A=> C(	1517	),
	B=>E(	1368	),
	Cin=> Carry( 	1452	),
	Cout=> Carry( 	1453	),
	S=> E(	1430	));
			
 U1454	: Somador_Exato_1 PORT MAP(
	A=> C(	1518	),
	B=>E(	1369	),
	Cin=> Carry( 	1453	),
	Cout=> Carry( 	1454	),
	S=> E(	1431	));
			
 U1455	: Somador_Exato_1 PORT MAP(
	A=> C(	1519	),
	B=>E(	1370	),
	Cin=> Carry( 	1454	),
	Cout=> Carry( 	1455	),
	S=> E(	1432	));
			
 U1456	: Somador_Exato_1 PORT MAP(
	A=> C(	1520	),
	B=>E(	1371	),
	Cin=> Carry( 	1455	),
	Cout=> Carry( 	1456	),
	S=> E(	1433	));
			
 U1457	: Somador_Exato_1 PORT MAP(
	A=> C(	1521	),
	B=>E(	1372	),
	Cin=> Carry( 	1456	),
	Cout=> Carry( 	1457	),
	S=> E(	1434	));
			
 U1458	: Somador_Exato_1 PORT MAP(
	A=> C(	1522	),
	B=>E(	1373	),
	Cin=> Carry( 	1457	),
	Cout=> Carry( 	1458	),
	S=> E(	1435	));
			
 U1459	: Somador_Exato_1 PORT MAP(
	A=> C(	1523	),
	B=>E(	1374	),
	Cin=> Carry( 	1458	),
	Cout=> Carry( 	1459	),
	S=> E(	1436	));
			
 U1460	: Somador_Exato_1 PORT MAP(
	A=> C(	1524	),
	B=>E(	1375	),
	Cin=> Carry( 	1459	),
	Cout=> Carry( 	1460	),
	S=> E(	1437	));
			
 U1461	: Somador_Exato_1 PORT MAP(
	A=> C(	1525	),
	B=>E(	1376	),
	Cin=> Carry( 	1460	),
	Cout=> Carry( 	1461	),
	S=> E(	1438	));
			
 U1462	: Somador_Exato_1 PORT MAP(
	A=> C(	1526	),
	B=>E(	1377	),
	Cin=> Carry( 	1461	),
	Cout=> Carry( 	1462	),
	S=> E(	1439	));
			
 U1463	: Somador_Exato_1 PORT MAP(
	A=> C(	1527	),
	B=>E(	1378	),
	Cin=> Carry( 	1462	),
	Cout=> Carry( 	1463	),
	S=> E(	1440	));
			
 U1464	: Somador_Exato_1 PORT MAP(
	A=> C(	1528	),
	B=>E(	1379	),
	Cin=> Carry( 	1463	),
	Cout=> Carry( 	1464	),
	S=> E(	1441	));
			
 U1465	: Somador_Exato_1 PORT MAP(
	A=> C(	1529	),
	B=>E(	1380	),
	Cin=> Carry( 	1464	),
	Cout=> Carry( 	1465	),
	S=> E(	1442	));
			
 U1466	: Somador_Exato_1 PORT MAP(
	A=> C(	1530	),
	B=>E(	1381	),
	Cin=> Carry( 	1465	),
	Cout=> Carry( 	1466	),
	S=> E(	1443	));
			
 U1467	: Somador_Exato_1 PORT MAP(
	A=> C(	1531	),
	B=>E(	1382	),
	Cin=> Carry( 	1466	),
	Cout=> Carry( 	1467	),
	S=> E(	1444	));
			
 U1468	: Somador_Exato_1 PORT MAP(
	A=> C(	1532	),
	B=>E(	1383	),
	Cin=> Carry( 	1467	),
	Cout=> Carry( 	1468	),
	S=> E(	1445	));
			
 U1469	: Somador_Exato_1 PORT MAP(
	A=> C(	1533	),
	B=>E(	1384	),
	Cin=> Carry( 	1468	),
	Cout=> Carry( 	1469	),
	S=> E(	1446	));
			
 U1470	: Somador_Exato_1 PORT MAP(
	A=> C(	1534	),
	B=>E(	1385	),
	Cin=> Carry( 	1469	),
	Cout=> Carry( 	1470	),
	S=> E(	1447	));
			
 U1471	: Somador_Exato_1 PORT MAP(
	A=> C(	1535	),
	B=>Carry(	1407	),
	Cin=> Carry( 	1470	),
	Cout=> Carry( 	1471	),
	S=> E(	1448	));

			
 U1472	: Somador_Exato_1 PORT MAP(
	A=> C(	1536	),
	B=>E(	1386	),
	Cin=> '0'	,
	Cout=> Carry( 	1472	),
	S=> R(	24	));
			
 U1473	: Somador_Exato_1 PORT MAP(
	A=> C(	1537	),
	B=>E(	1387	),
	Cin=> Carry( 	1472	),
	Cout=> Carry( 	1473	),
	S=> E(	1449	));
			
 U1474	: Somador_Exato_1 PORT MAP(
	A=> C(	1538	),
	B=>E(	1388	),
	Cin=> Carry( 	1473	),
	Cout=> Carry( 	1474	),
	S=> E(	1450	));
			
 U1475	: Somador_Exato_1 PORT MAP(
	A=> C(	1539	),
	B=>E(	1389	),
	Cin=> Carry( 	1474	),
	Cout=> Carry( 	1475	),
	S=> E(	1451	));
			
 U1476	: Somador_Exato_1 PORT MAP(
	A=> C(	1540	),
	B=>E(	1390	),
	Cin=> Carry( 	1475	),
	Cout=> Carry( 	1476	),
	S=> E(	1452	));
			
 U1477	: Somador_Exato_1 PORT MAP(
	A=> C(	1541	),
	B=>E(	1391	),
	Cin=> Carry( 	1476	),
	Cout=> Carry( 	1477	),
	S=> E(	1453	));
			
 U1478	: Somador_Exato_1 PORT MAP(
	A=> C(	1542	),
	B=>E(	1392	),
	Cin=> Carry( 	1477	),
	Cout=> Carry( 	1478	),
	S=> E(	1454	));
			
 U1479	: Somador_Exato_1 PORT MAP(
	A=> C(	1543	),
	B=>E(	1393	),
	Cin=> Carry( 	1478	),
	Cout=> Carry( 	1479	),
	S=> E(	1455	));
			
 U1480	: Somador_Exato_1 PORT MAP(
	A=> C(	1544	),
	B=>E(	1394	),
	Cin=> Carry( 	1479	),
	Cout=> Carry( 	1480	),
	S=> E(	1456	));
			
 U1481	: Somador_Exato_1 PORT MAP(
	A=> C(	1545	),
	B=>E(	1395	),
	Cin=> Carry( 	1480	),
	Cout=> Carry( 	1481	),
	S=> E(	1457	));
			
 U1482	: Somador_Exato_1 PORT MAP(
	A=> C(	1546	),
	B=>E(	1396	),
	Cin=> Carry( 	1481	),
	Cout=> Carry( 	1482	),
	S=> E(	1458	));
			
 U1483	: Somador_Exato_1 PORT MAP(
	A=> C(	1547	),
	B=>E(	1397	),
	Cin=> Carry( 	1482	),
	Cout=> Carry( 	1483	),
	S=> E(	1459	));
			
 U1484	: Somador_Exato_1 PORT MAP(
	A=> C(	1548	),
	B=>E(	1398	),
	Cin=> Carry( 	1483	),
	Cout=> Carry( 	1484	),
	S=> E(	1460	));
			
 U1485	: Somador_Exato_1 PORT MAP(
	A=> C(	1549	),
	B=>E(	1399	),
	Cin=> Carry( 	1484	),
	Cout=> Carry( 	1485	),
	S=> E(	1461	));
			
 U1486	: Somador_Exato_1 PORT MAP(
	A=> C(	1550	),
	B=>E(	1400	),
	Cin=> Carry( 	1485	),
	Cout=> Carry( 	1486	),
	S=> E(	1462	));
			
 U1487	: Somador_Exato_1 PORT MAP(
	A=> C(	1551	),
	B=>E(	1401	),
	Cin=> Carry( 	1486	),
	Cout=> Carry( 	1487	),
	S=> E(	1463	));
			
 U1488	: Somador_Exato_1 PORT MAP(
	A=> C(	1552	),
	B=>E(	1402	),
	Cin=> Carry( 	1487	),
	Cout=> Carry( 	1488	),
	S=> E(	1464	));
			
 U1489	: Somador_Exato_1 PORT MAP(
	A=> C(	1553	),
	B=>E(	1403	),
	Cin=> Carry( 	1488	),
	Cout=> Carry( 	1489	),
	S=> E(	1465	));
			
 U1490	: Somador_Exato_1 PORT MAP(
	A=> C(	1554	),
	B=>E(	1404	),
	Cin=> Carry( 	1489	),
	Cout=> Carry( 	1490	),
	S=> E(	1466	));
			
 U1491	: Somador_Exato_1 PORT MAP(
	A=> C(	1555	),
	B=>E(	1405	),
	Cin=> Carry( 	1490	),
	Cout=> Carry( 	1491	),
	S=> E(	1467	));
			
 U1492	: Somador_Exato_1 PORT MAP(
	A=> C(	1556	),
	B=>E(	1406	),
	Cin=> Carry( 	1491	),
	Cout=> Carry( 	1492	),
	S=> E(	1468	));
			
 U1493	: Somador_Exato_1 PORT MAP(
	A=> C(	1557	),
	B=>E(	1407	),
	Cin=> Carry( 	1492	),
	Cout=> Carry( 	1493	),
	S=> E(	1469	));
			
 U1494	: Somador_Exato_1 PORT MAP(
	A=> C(	1558	),
	B=>E(	1408	),
	Cin=> Carry( 	1493	),
	Cout=> Carry( 	1494	),
	S=> E(	1470	));
			
 U1495	: Somador_Exato_1 PORT MAP(
	A=> C(	1559	),
	B=>E(	1409	),
	Cin=> Carry( 	1494	),
	Cout=> Carry( 	1495	),
	S=> E(	1471	));
			
 U1496	: Somador_Exato_1 PORT MAP(
	A=> C(	1560	),
	B=>E(	1410	),
	Cin=> Carry( 	1495	),
	Cout=> Carry( 	1496	),
	S=> E(	1472	));
			
 U1497	: Somador_Exato_1 PORT MAP(
	A=> C(	1561	),
	B=>E(	1411	),
	Cin=> Carry( 	1496	),
	Cout=> Carry( 	1497	),
	S=> E(	1473	));
			
 U1498	: Somador_Exato_1 PORT MAP(
	A=> C(	1562	),
	B=>E(	1412	),
	Cin=> Carry( 	1497	),
	Cout=> Carry( 	1498	),
	S=> E(	1474	));
			
 U1499	: Somador_Exato_1 PORT MAP(
	A=> C(	1563	),
	B=>E(	1413	),
	Cin=> Carry( 	1498	),
	Cout=> Carry( 	1499	),
	S=> E(	1475	));
			
 U1500	: Somador_Exato_1 PORT MAP(
	A=> C(	1564	),
	B=>E(	1414	),
	Cin=> Carry( 	1499	),
	Cout=> Carry( 	1500	),
	S=> E(	1476	));
			
 U1501	: Somador_Exato_1 PORT MAP(
	A=> C(	1565	),
	B=>E(	1415	),
	Cin=> Carry( 	1500	),
	Cout=> Carry( 	1501	),
	S=> E(	1477	));
			
 U1502	: Somador_Exato_1 PORT MAP(
	A=> C(	1566	),
	B=>E(	1416	),
	Cin=> Carry( 	1501	),
	Cout=> Carry( 	1502	),
	S=> E(	1478	));
			
 U1503	: Somador_Exato_1 PORT MAP(
	A=> C(	1567	),
	B=>E(	1417	),
	Cin=> Carry( 	1502	),
	Cout=> Carry( 	1503	),
	S=> E(	1479	));
			
 U1504	: Somador_Exato_1 PORT MAP(
	A=> C(	1568	),
	B=>E(	1418	),
	Cin=> Carry( 	1503	),
	Cout=> Carry( 	1504	),
	S=> E(	1480	));
			
 U1505	: Somador_Exato_1 PORT MAP(
	A=> C(	1569	),
	B=>E(	1419	),
	Cin=> Carry( 	1504	),
	Cout=> Carry( 	1505	),
	S=> E(	1481	));
			
 U1506	: Somador_Exato_1 PORT MAP(
	A=> C(	1570	),
	B=>E(	1420	),
	Cin=> Carry( 	1505	),
	Cout=> Carry( 	1506	),
	S=> E(	1482	));
			
 U1507	: Somador_Exato_1 PORT MAP(
	A=> C(	1571	),
	B=>E(	1421	),
	Cin=> Carry( 	1506	),
	Cout=> Carry( 	1507	),
	S=> E(	1483	));
			
 U1508	: Somador_Exato_1 PORT MAP(
	A=> C(	1572	),
	B=>E(	1422	),
	Cin=> Carry( 	1507	),
	Cout=> Carry( 	1508	),
	S=> E(	1484	));
			
 U1509	: Somador_Exato_1 PORT MAP(
	A=> C(	1573	),
	B=>E(	1423	),
	Cin=> Carry( 	1508	),
	Cout=> Carry( 	1509	),
	S=> E(	1485	));
			
 U1510	: Somador_Exato_1 PORT MAP(
	A=> C(	1574	),
	B=>E(	1424	),
	Cin=> Carry( 	1509	),
	Cout=> Carry( 	1510	),
	S=> E(	1486	));
			
 U1511	: Somador_Exato_1 PORT MAP(
	A=> C(	1575	),
	B=>E(	1425	),
	Cin=> Carry( 	1510	),
	Cout=> Carry( 	1511	),
	S=> E(	1487	));
			
 U1512	: Somador_Exato_1 PORT MAP(
	A=> C(	1576	),
	B=>E(	1426	),
	Cin=> Carry( 	1511	),
	Cout=> Carry( 	1512	),
	S=> E(	1488	));
			
 U1513	: Somador_Exato_1 PORT MAP(
	A=> C(	1577	),
	B=>E(	1427	),
	Cin=> Carry( 	1512	),
	Cout=> Carry( 	1513	),
	S=> E(	1489	));
			
 U1514	: Somador_Exato_1 PORT MAP(
	A=> C(	1578	),
	B=>E(	1428	),
	Cin=> Carry( 	1513	),
	Cout=> Carry( 	1514	),
	S=> E(	1490	));
			
 U1515	: Somador_Exato_1 PORT MAP(
	A=> C(	1579	),
	B=>E(	1429	),
	Cin=> Carry( 	1514	),
	Cout=> Carry( 	1515	),
	S=> E(	1491	));
			
 U1516	: Somador_Exato_1 PORT MAP(
	A=> C(	1580	),
	B=>E(	1430	),
	Cin=> Carry( 	1515	),
	Cout=> Carry( 	1516	),
	S=> E(	1492	));
			
 U1517	: Somador_Exato_1 PORT MAP(
	A=> C(	1581	),
	B=>E(	1431	),
	Cin=> Carry( 	1516	),
	Cout=> Carry( 	1517	),
	S=> E(	1493	));
			
 U1518	: Somador_Exato_1 PORT MAP(
	A=> C(	1582	),
	B=>E(	1432	),
	Cin=> Carry( 	1517	),
	Cout=> Carry( 	1518	),
	S=> E(	1494	));
			
 U1519	: Somador_Exato_1 PORT MAP(
	A=> C(	1583	),
	B=>E(	1433	),
	Cin=> Carry( 	1518	),
	Cout=> Carry( 	1519	),
	S=> E(	1495	));
			
 U1520	: Somador_Exato_1 PORT MAP(
	A=> C(	1584	),
	B=>E(	1434	),
	Cin=> Carry( 	1519	),
	Cout=> Carry( 	1520	),
	S=> E(	1496	));
			
 U1521	: Somador_Exato_1 PORT MAP(
	A=> C(	1585	),
	B=>E(	1435	),
	Cin=> Carry( 	1520	),
	Cout=> Carry( 	1521	),
	S=> E(	1497	));
			
 U1522	: Somador_Exato_1 PORT MAP(
	A=> C(	1586	),
	B=>E(	1436	),
	Cin=> Carry( 	1521	),
	Cout=> Carry( 	1522	),
	S=> E(	1498	));
			
 U1523	: Somador_Exato_1 PORT MAP(
	A=> C(	1587	),
	B=>E(	1437	),
	Cin=> Carry( 	1522	),
	Cout=> Carry( 	1523	),
	S=> E(	1499	));
			
 U1524	: Somador_Exato_1 PORT MAP(
	A=> C(	1588	),
	B=>E(	1438	),
	Cin=> Carry( 	1523	),
	Cout=> Carry( 	1524	),
	S=> E(	1500	));
			
 U1525	: Somador_Exato_1 PORT MAP(
	A=> C(	1589	),
	B=>E(	1439	),
	Cin=> Carry( 	1524	),
	Cout=> Carry( 	1525	),
	S=> E(	1501	));
			
 U1526	: Somador_Exato_1 PORT MAP(
	A=> C(	1590	),
	B=>E(	1440	),
	Cin=> Carry( 	1525	),
	Cout=> Carry( 	1526	),
	S=> E(	1502	));
			
 U1527	: Somador_Exato_1 PORT MAP(
	A=> C(	1591	),
	B=>E(	1441	),
	Cin=> Carry( 	1526	),
	Cout=> Carry( 	1527	),
	S=> E(	1503	));
			
 U1528	: Somador_Exato_1 PORT MAP(
	A=> C(	1592	),
	B=>E(	1442	),
	Cin=> Carry( 	1527	),
	Cout=> Carry( 	1528	),
	S=> E(	1504	));
			
 U1529	: Somador_Exato_1 PORT MAP(
	A=> C(	1593	),
	B=>E(	1443	),
	Cin=> Carry( 	1528	),
	Cout=> Carry( 	1529	),
	S=> E(	1505	));
			
 U1530	: Somador_Exato_1 PORT MAP(
	A=> C(	1594	),
	B=>E(	1444	),
	Cin=> Carry( 	1529	),
	Cout=> Carry( 	1530	),
	S=> E(	1506	));
			
 U1531	: Somador_Exato_1 PORT MAP(
	A=> C(	1595	),
	B=>E(	1445	),
	Cin=> Carry( 	1530	),
	Cout=> Carry( 	1531	),
	S=> E(	1507	));
			
 U1532	: Somador_Exato_1 PORT MAP(
	A=> C(	1596	),
	B=>E(	1446	),
	Cin=> Carry( 	1531	),
	Cout=> Carry( 	1532	),
	S=> E(	1508	));
			
 U1533	: Somador_Exato_1 PORT MAP(
	A=> C(	1597	),
	B=>E(	1447	),
	Cin=> Carry( 	1532	),
	Cout=> Carry( 	1533	),
	S=> E(	1509	));
			
 U1534	: Somador_Exato_1 PORT MAP(
	A=> C(	1598	),
	B=>E(	1448	),
	Cin=> Carry( 	1533	),
	Cout=> Carry( 	1534	),
	S=> E(	1510	));
			
 U1535	: Somador_Exato_1 PORT MAP(
	A=> C(	1599	),
	B=>Carry(	1471	),
	Cin=> Carry( 	1534	),
	Cout=> Carry( 	1535	),
	S=> E(	1511	));

			
 U1536	: Somador_Exato_1 PORT MAP(
	A=> C(	1600	),
	B=>E(	1449	),
	Cin=> '0'	,
	Cout=> Carry( 	1536	),
	S=> R(	25	));
			
 U1537	: Somador_Exato_1 PORT MAP(
	A=> C(	1601	),
	B=>E(	1450	),
	Cin=> Carry( 	1536	),
	Cout=> Carry( 	1537	),
	S=> E(	1512	));
			
 U1538	: Somador_Exato_1 PORT MAP(
	A=> C(	1602	),
	B=>E(	1451	),
	Cin=> Carry( 	1537	),
	Cout=> Carry( 	1538	),
	S=> E(	1513	));
			
 U1539	: Somador_Exato_1 PORT MAP(
	A=> C(	1603	),
	B=>E(	1452	),
	Cin=> Carry( 	1538	),
	Cout=> Carry( 	1539	),
	S=> E(	1514	));
			
 U1540	: Somador_Exato_1 PORT MAP(
	A=> C(	1604	),
	B=>E(	1453	),
	Cin=> Carry( 	1539	),
	Cout=> Carry( 	1540	),
	S=> E(	1515	));
			
 U1541	: Somador_Exato_1 PORT MAP(
	A=> C(	1605	),
	B=>E(	1454	),
	Cin=> Carry( 	1540	),
	Cout=> Carry( 	1541	),
	S=> E(	1516	));
			
 U1542	: Somador_Exato_1 PORT MAP(
	A=> C(	1606	),
	B=>E(	1455	),
	Cin=> Carry( 	1541	),
	Cout=> Carry( 	1542	),
	S=> E(	1517	));
			
 U1543	: Somador_Exato_1 PORT MAP(
	A=> C(	1607	),
	B=>E(	1456	),
	Cin=> Carry( 	1542	),
	Cout=> Carry( 	1543	),
	S=> E(	1518	));
			
 U1544	: Somador_Exato_1 PORT MAP(
	A=> C(	1608	),
	B=>E(	1457	),
	Cin=> Carry( 	1543	),
	Cout=> Carry( 	1544	),
	S=> E(	1519	));
			
 U1545	: Somador_Exato_1 PORT MAP(
	A=> C(	1609	),
	B=>E(	1458	),
	Cin=> Carry( 	1544	),
	Cout=> Carry( 	1545	),
	S=> E(	1520	));
			
 U1546	: Somador_Exato_1 PORT MAP(
	A=> C(	1610	),
	B=>E(	1459	),
	Cin=> Carry( 	1545	),
	Cout=> Carry( 	1546	),
	S=> E(	1521	));
			
 U1547	: Somador_Exato_1 PORT MAP(
	A=> C(	1611	),
	B=>E(	1460	),
	Cin=> Carry( 	1546	),
	Cout=> Carry( 	1547	),
	S=> E(	1522	));
			
 U1548	: Somador_Exato_1 PORT MAP(
	A=> C(	1612	),
	B=>E(	1461	),
	Cin=> Carry( 	1547	),
	Cout=> Carry( 	1548	),
	S=> E(	1523	));
			
 U1549	: Somador_Exato_1 PORT MAP(
	A=> C(	1613	),
	B=>E(	1462	),
	Cin=> Carry( 	1548	),
	Cout=> Carry( 	1549	),
	S=> E(	1524	));
			
 U1550	: Somador_Exato_1 PORT MAP(
	A=> C(	1614	),
	B=>E(	1463	),
	Cin=> Carry( 	1549	),
	Cout=> Carry( 	1550	),
	S=> E(	1525	));
			
 U1551	: Somador_Exato_1 PORT MAP(
	A=> C(	1615	),
	B=>E(	1464	),
	Cin=> Carry( 	1550	),
	Cout=> Carry( 	1551	),
	S=> E(	1526	));
			
 U1552	: Somador_Exato_1 PORT MAP(
	A=> C(	1616	),
	B=>E(	1465	),
	Cin=> Carry( 	1551	),
	Cout=> Carry( 	1552	),
	S=> E(	1527	));
			
 U1553	: Somador_Exato_1 PORT MAP(
	A=> C(	1617	),
	B=>E(	1466	),
	Cin=> Carry( 	1552	),
	Cout=> Carry( 	1553	),
	S=> E(	1528	));
			
 U1554	: Somador_Exato_1 PORT MAP(
	A=> C(	1618	),
	B=>E(	1467	),
	Cin=> Carry( 	1553	),
	Cout=> Carry( 	1554	),
	S=> E(	1529	));
			
 U1555	: Somador_Exato_1 PORT MAP(
	A=> C(	1619	),
	B=>E(	1468	),
	Cin=> Carry( 	1554	),
	Cout=> Carry( 	1555	),
	S=> E(	1530	));
			
 U1556	: Somador_Exato_1 PORT MAP(
	A=> C(	1620	),
	B=>E(	1469	),
	Cin=> Carry( 	1555	),
	Cout=> Carry( 	1556	),
	S=> E(	1531	));
			
 U1557	: Somador_Exato_1 PORT MAP(
	A=> C(	1621	),
	B=>E(	1470	),
	Cin=> Carry( 	1556	),
	Cout=> Carry( 	1557	),
	S=> E(	1532	));
			
 U1558	: Somador_Exato_1 PORT MAP(
	A=> C(	1622	),
	B=>E(	1471	),
	Cin=> Carry( 	1557	),
	Cout=> Carry( 	1558	),
	S=> E(	1533	));
			
 U1559	: Somador_Exato_1 PORT MAP(
	A=> C(	1623	),
	B=>E(	1472	),
	Cin=> Carry( 	1558	),
	Cout=> Carry( 	1559	),
	S=> E(	1534	));
			
 U1560	: Somador_Exato_1 PORT MAP(
	A=> C(	1624	),
	B=>E(	1473	),
	Cin=> Carry( 	1559	),
	Cout=> Carry( 	1560	),
	S=> E(	1535	));
			
 U1561	: Somador_Exato_1 PORT MAP(
	A=> C(	1625	),
	B=>E(	1474	),
	Cin=> Carry( 	1560	),
	Cout=> Carry( 	1561	),
	S=> E(	1536	));
			
 U1562	: Somador_Exato_1 PORT MAP(
	A=> C(	1626	),
	B=>E(	1475	),
	Cin=> Carry( 	1561	),
	Cout=> Carry( 	1562	),
	S=> E(	1537	));
			
 U1563	: Somador_Exato_1 PORT MAP(
	A=> C(	1627	),
	B=>E(	1476	),
	Cin=> Carry( 	1562	),
	Cout=> Carry( 	1563	),
	S=> E(	1538	));
			
 U1564	: Somador_Exato_1 PORT MAP(
	A=> C(	1628	),
	B=>E(	1477	),
	Cin=> Carry( 	1563	),
	Cout=> Carry( 	1564	),
	S=> E(	1539	));
			
 U1565	: Somador_Exato_1 PORT MAP(
	A=> C(	1629	),
	B=>E(	1478	),
	Cin=> Carry( 	1564	),
	Cout=> Carry( 	1565	),
	S=> E(	1540	));
			
 U1566	: Somador_Exato_1 PORT MAP(
	A=> C(	1630	),
	B=>E(	1479	),
	Cin=> Carry( 	1565	),
	Cout=> Carry( 	1566	),
	S=> E(	1541	));
			
 U1567	: Somador_Exato_1 PORT MAP(
	A=> C(	1631	),
	B=>E(	1480	),
	Cin=> Carry( 	1566	),
	Cout=> Carry( 	1567	),
	S=> E(	1542	));
			
 U1568	: Somador_Exato_1 PORT MAP(
	A=> C(	1632	),
	B=>E(	1481	),
	Cin=> Carry( 	1567	),
	Cout=> Carry( 	1568	),
	S=> E(	1543	));
			
 U1569	: Somador_Exato_1 PORT MAP(
	A=> C(	1633	),
	B=>E(	1482	),
	Cin=> Carry( 	1568	),
	Cout=> Carry( 	1569	),
	S=> E(	1544	));
			
 U1570	: Somador_Exato_1 PORT MAP(
	A=> C(	1634	),
	B=>E(	1483	),
	Cin=> Carry( 	1569	),
	Cout=> Carry( 	1570	),
	S=> E(	1545	));
			
 U1571	: Somador_Exato_1 PORT MAP(
	A=> C(	1635	),
	B=>E(	1484	),
	Cin=> Carry( 	1570	),
	Cout=> Carry( 	1571	),
	S=> E(	1546	));
			
 U1572	: Somador_Exato_1 PORT MAP(
	A=> C(	1636	),
	B=>E(	1485	),
	Cin=> Carry( 	1571	),
	Cout=> Carry( 	1572	),
	S=> E(	1547	));
			
 U1573	: Somador_Exato_1 PORT MAP(
	A=> C(	1637	),
	B=>E(	1486	),
	Cin=> Carry( 	1572	),
	Cout=> Carry( 	1573	),
	S=> E(	1548	));
			
 U1574	: Somador_Exato_1 PORT MAP(
	A=> C(	1638	),
	B=>E(	1487	),
	Cin=> Carry( 	1573	),
	Cout=> Carry( 	1574	),
	S=> E(	1549	));
			
 U1575	: Somador_Exato_1 PORT MAP(
	A=> C(	1639	),
	B=>E(	1488	),
	Cin=> Carry( 	1574	),
	Cout=> Carry( 	1575	),
	S=> E(	1550	));
			
 U1576	: Somador_Exato_1 PORT MAP(
	A=> C(	1640	),
	B=>E(	1489	),
	Cin=> Carry( 	1575	),
	Cout=> Carry( 	1576	),
	S=> E(	1551	));
			
 U1577	: Somador_Exato_1 PORT MAP(
	A=> C(	1641	),
	B=>E(	1490	),
	Cin=> Carry( 	1576	),
	Cout=> Carry( 	1577	),
	S=> E(	1552	));
			
 U1578	: Somador_Exato_1 PORT MAP(
	A=> C(	1642	),
	B=>E(	1491	),
	Cin=> Carry( 	1577	),
	Cout=> Carry( 	1578	),
	S=> E(	1553	));
			
 U1579	: Somador_Exato_1 PORT MAP(
	A=> C(	1643	),
	B=>E(	1492	),
	Cin=> Carry( 	1578	),
	Cout=> Carry( 	1579	),
	S=> E(	1554	));
			
 U1580	: Somador_Exato_1 PORT MAP(
	A=> C(	1644	),
	B=>E(	1493	),
	Cin=> Carry( 	1579	),
	Cout=> Carry( 	1580	),
	S=> E(	1555	));
			
 U1581	: Somador_Exato_1 PORT MAP(
	A=> C(	1645	),
	B=>E(	1494	),
	Cin=> Carry( 	1580	),
	Cout=> Carry( 	1581	),
	S=> E(	1556	));
			
 U1582	: Somador_Exato_1 PORT MAP(
	A=> C(	1646	),
	B=>E(	1495	),
	Cin=> Carry( 	1581	),
	Cout=> Carry( 	1582	),
	S=> E(	1557	));
			
 U1583	: Somador_Exato_1 PORT MAP(
	A=> C(	1647	),
	B=>E(	1496	),
	Cin=> Carry( 	1582	),
	Cout=> Carry( 	1583	),
	S=> E(	1558	));
			
 U1584	: Somador_Exato_1 PORT MAP(
	A=> C(	1648	),
	B=>E(	1497	),
	Cin=> Carry( 	1583	),
	Cout=> Carry( 	1584	),
	S=> E(	1559	));
			
 U1585	: Somador_Exato_1 PORT MAP(
	A=> C(	1649	),
	B=>E(	1498	),
	Cin=> Carry( 	1584	),
	Cout=> Carry( 	1585	),
	S=> E(	1560	));
			
 U1586	: Somador_Exato_1 PORT MAP(
	A=> C(	1650	),
	B=>E(	1499	),
	Cin=> Carry( 	1585	),
	Cout=> Carry( 	1586	),
	S=> E(	1561	));
			
 U1587	: Somador_Exato_1 PORT MAP(
	A=> C(	1651	),
	B=>E(	1500	),
	Cin=> Carry( 	1586	),
	Cout=> Carry( 	1587	),
	S=> E(	1562	));
			
 U1588	: Somador_Exato_1 PORT MAP(
	A=> C(	1652	),
	B=>E(	1501	),
	Cin=> Carry( 	1587	),
	Cout=> Carry( 	1588	),
	S=> E(	1563	));
			
 U1589	: Somador_Exato_1 PORT MAP(
	A=> C(	1653	),
	B=>E(	1502	),
	Cin=> Carry( 	1588	),
	Cout=> Carry( 	1589	),
	S=> E(	1564	));
			
 U1590	: Somador_Exato_1 PORT MAP(
	A=> C(	1654	),
	B=>E(	1503	),
	Cin=> Carry( 	1589	),
	Cout=> Carry( 	1590	),
	S=> E(	1565	));
			
 U1591	: Somador_Exato_1 PORT MAP(
	A=> C(	1655	),
	B=>E(	1504	),
	Cin=> Carry( 	1590	),
	Cout=> Carry( 	1591	),
	S=> E(	1566	));
			
 U1592	: Somador_Exato_1 PORT MAP(
	A=> C(	1656	),
	B=>E(	1505	),
	Cin=> Carry( 	1591	),
	Cout=> Carry( 	1592	),
	S=> E(	1567	));
			
 U1593	: Somador_Exato_1 PORT MAP(
	A=> C(	1657	),
	B=>E(	1506	),
	Cin=> Carry( 	1592	),
	Cout=> Carry( 	1593	),
	S=> E(	1568	));
			
 U1594	: Somador_Exato_1 PORT MAP(
	A=> C(	1658	),
	B=>E(	1507	),
	Cin=> Carry( 	1593	),
	Cout=> Carry( 	1594	),
	S=> E(	1569	));
			
 U1595	: Somador_Exato_1 PORT MAP(
	A=> C(	1659	),
	B=>E(	1508	),
	Cin=> Carry( 	1594	),
	Cout=> Carry( 	1595	),
	S=> E(	1570	));
			
 U1596	: Somador_Exato_1 PORT MAP(
	A=> C(	1660	),
	B=>E(	1509	),
	Cin=> Carry( 	1595	),
	Cout=> Carry( 	1596	),
	S=> E(	1571	));
			
 U1597	: Somador_Exato_1 PORT MAP(
	A=> C(	1661	),
	B=>E(	1510	),
	Cin=> Carry( 	1596	),
	Cout=> Carry( 	1597	),
	S=> E(	1572	));
			
 U1598	: Somador_Exato_1 PORT MAP(
	A=> C(	1662	),
	B=>E(	1511	),
	Cin=> Carry( 	1597	),
	Cout=> Carry( 	1598	),
	S=> E(	1573	));
			
 U1599	: Somador_Exato_1 PORT MAP(
	A=> C(	1663	),
	B=>Carry(	1535	),
	Cin=> Carry( 	1598	),
	Cout=> Carry( 	1599	),
	S=> E(	1574	));

			
 U1600	: Somador_Exato_1 PORT MAP(
	A=> C(	1664	),
	B=>E(	1512	),
	Cin=> '0'	,
	Cout=> Carry( 	1600	),
	S=> R(	26	));
			
  U1601	: Somador_Exato_1 PORT MAP(
	A=> C(	1665	),
	B=>E(	1513	),
	Cin=> Carry( 	1600	),
	Cout=> Carry( 	1601	),
	S=> E(	1575	));
			
  U1602	: Somador_Exato_1 PORT MAP(
	A=> C(	1666	),
	B=>E(	1514	),
	Cin=> Carry( 	1601	),
	Cout=> Carry( 	1602	),
	S=> E(	1576	));
			
  U1603	: Somador_Exato_1 PORT MAP(
	A=> C(	1667	),
	B=>E(	1515	),
	Cin=> Carry( 	1602	),
	Cout=> Carry( 	1603	),
	S=> E(	1577	));
			
  U1604	: Somador_Exato_1 PORT MAP(
	A=> C(	1668	),
	B=>E(	1516	),
	Cin=> Carry( 	1603	),
	Cout=> Carry( 	1604	),
	S=> E(	1578	));
			
  U1605	: Somador_Exato_1 PORT MAP(
	A=> C(	1669	),
	B=>E(	1517	),
	Cin=> Carry( 	1604	),
	Cout=> Carry( 	1605	),
	S=> E(	1579	));
			
  U1606	: Somador_Exato_1 PORT MAP(
	A=> C(	1670	),
	B=>E(	1518	),
	Cin=> Carry( 	1605	),
	Cout=> Carry( 	1606	),
	S=> E(	1580	));
			
  U1607	: Somador_Exato_1 PORT MAP(
	A=> C(	1671	),
	B=>E(	1519	),
	Cin=> Carry( 	1606	),
	Cout=> Carry( 	1607	),
	S=> E(	1581	));
			
  U1608	: Somador_Exato_1 PORT MAP(
	A=> C(	1672	),
	B=>E(	1520	),
	Cin=> Carry( 	1607	),
	Cout=> Carry( 	1608	),
	S=> E(	1582	));
			
  U1609	: Somador_Exato_1 PORT MAP(
	A=> C(	1673	),
	B=>E(	1521	),
	Cin=> Carry( 	1608	),
	Cout=> Carry( 	1609	),
	S=> E(	1583	));
			
  U1610	: Somador_Exato_1 PORT MAP(
	A=> C(	1674	),
	B=>E(	1522	),
	Cin=> Carry( 	1609	),
	Cout=> Carry( 	1610	),
	S=> E(	1584	));
			
  U1611	: Somador_Exato_1 PORT MAP(
	A=> C(	1675	),
	B=>E(	1523	),
	Cin=> Carry( 	1610	),
	Cout=> Carry( 	1611	),
	S=> E(	1585	));
			
  U1612	: Somador_Exato_1 PORT MAP(
	A=> C(	1676	),
	B=>E(	1524	),
	Cin=> Carry( 	1611	),
	Cout=> Carry( 	1612	),
	S=> E(	1586	));
			
  U1613	: Somador_Exato_1 PORT MAP(
	A=> C(	1677	),
	B=>E(	1525	),
	Cin=> Carry( 	1612	),
	Cout=> Carry( 	1613	),
	S=> E(	1587	));
			
  U1614	: Somador_Exato_1 PORT MAP(
	A=> C(	1678	),
	B=>E(	1526	),
	Cin=> Carry( 	1613	),
	Cout=> Carry( 	1614	),
	S=> E(	1588	));
			
  U1615	: Somador_Exato_1 PORT MAP(
	A=> C(	1679	),
	B=>E(	1527	),
	Cin=> Carry( 	1614	),
	Cout=> Carry( 	1615	),
	S=> E(	1589	));
			
  U1616	: Somador_Exato_1 PORT MAP(
	A=> C(	1680	),
	B=>E(	1528	),
	Cin=> Carry( 	1615	),
	Cout=> Carry( 	1616	),
	S=> E(	1590	));
			
  U1617	: Somador_Exato_1 PORT MAP(
	A=> C(	1681	),
	B=>E(	1529	),
	Cin=> Carry( 	1616	),
	Cout=> Carry( 	1617	),
	S=> E(	1591	));
			
  U1618	: Somador_Exato_1 PORT MAP(
	A=> C(	1682	),
	B=>E(	1530	),
	Cin=> Carry( 	1617	),
	Cout=> Carry( 	1618	),
	S=> E(	1592	));
			
  U1619	: Somador_Exato_1 PORT MAP(
	A=> C(	1683	),
	B=>E(	1531	),
	Cin=> Carry( 	1618	),
	Cout=> Carry( 	1619	),
	S=> E(	1593	));
			
  U1620	: Somador_Exato_1 PORT MAP(
	A=> C(	1684	),
	B=>E(	1532	),
	Cin=> Carry( 	1619	),
	Cout=> Carry( 	1620	),
	S=> E(	1594	));
			
  U1621	: Somador_Exato_1 PORT MAP(
	A=> C(	1685	),
	B=>E(	1533	),
	Cin=> Carry( 	1620	),
	Cout=> Carry( 	1621	),
	S=> E(	1595	));
			
  U1622	: Somador_Exato_1 PORT MAP(
	A=> C(	1686	),
	B=>E(	1534	),
	Cin=> Carry( 	1621	),
	Cout=> Carry( 	1622	),
	S=> E(	1596	));
			
  U1623	: Somador_Exato_1 PORT MAP(
	A=> C(	1687	),
	B=>E(	1535	),
	Cin=> Carry( 	1622	),
	Cout=> Carry( 	1623	),
	S=> E(	1597	));
			
  U1624	: Somador_Exato_1 PORT MAP(
	A=> C(	1688	),
	B=>E(	1536	),
	Cin=> Carry( 	1623	),
	Cout=> Carry( 	1624	),
	S=> E(	1598	));
			
  U1625	: Somador_Exato_1 PORT MAP(
	A=> C(	1689	),
	B=>E(	1537	),
	Cin=> Carry( 	1624	),
	Cout=> Carry( 	1625	),
	S=> E(	1599	));
			
  U1626	: Somador_Exato_1 PORT MAP(
	A=> C(	1690	),
	B=>E(	1538	),
	Cin=> Carry( 	1625	),
	Cout=> Carry( 	1626	),
	S=> E(	1600	));
			
  U1627	: Somador_Exato_1 PORT MAP(
	A=> C(	1691	),
	B=>E(	1539	),
	Cin=> Carry( 	1626	),
	Cout=> Carry( 	1627	),
	S=> E(	1601	));
			
  U1628	: Somador_Exato_1 PORT MAP(
	A=> C(	1692	),
	B=>E(	1540	),
	Cin=> Carry( 	1627	),
	Cout=> Carry( 	1628	),
	S=> E(	1602	));
			
  U1629	: Somador_Exato_1 PORT MAP(
	A=> C(	1693	),
	B=>E(	1541	),
	Cin=> Carry( 	1628	),
	Cout=> Carry( 	1629	),
	S=> E(	1603	));
			
  U1630	: Somador_Exato_1 PORT MAP(
	A=> C(	1694	),
	B=>E(	1542	),
	Cin=> Carry( 	1629	),
	Cout=> Carry( 	1630	),
	S=> E(	1604	));
			
  U1631	: Somador_Exato_1 PORT MAP(
	A=> C(	1695	),
	B=>E(	1543	),
	Cin=> Carry( 	1630	),
	Cout=> Carry( 	1631	),
	S=> E(	1605	));
			
  U1632	: Somador_Exato_1 PORT MAP(
	A=> C(	1696	),
	B=>E(	1544	),
	Cin=> Carry( 	1631	),
	Cout=> Carry( 	1632	),
	S=> E(	1606	));
			
  U1633	: Somador_Exato_1 PORT MAP(
	A=> C(	1697	),
	B=>E(	1545	),
	Cin=> Carry( 	1632	),
	Cout=> Carry( 	1633	),
	S=> E(	1607	));
			
  U1634	: Somador_Exato_1 PORT MAP(
	A=> C(	1698	),
	B=>E(	1546	),
	Cin=> Carry( 	1633	),
	Cout=> Carry( 	1634	),
	S=> E(	1608	));
			
  U1635	: Somador_Exato_1 PORT MAP(
	A=> C(	1699	),
	B=>E(	1547	),
	Cin=> Carry( 	1634	),
	Cout=> Carry( 	1635	),
	S=> E(	1609	));
			
  U1636	: Somador_Exato_1 PORT MAP(
	A=> C(	1700	),
	B=>E(	1548	),
	Cin=> Carry( 	1635	),
	Cout=> Carry( 	1636	),
	S=> E(	1610	));
			
  U1637	: Somador_Exato_1 PORT MAP(
	A=> C(	1701	),
	B=>E(	1549	),
	Cin=> Carry( 	1636	),
	Cout=> Carry( 	1637	),
	S=> E(	1611	));
			
  U1638	: Somador_Exato_1 PORT MAP(
	A=> C(	1702	),
	B=>E(	1550	),
	Cin=> Carry( 	1637	),
	Cout=> Carry( 	1638	),
	S=> E(	1612	));
			
  U1639	: Somador_Exato_1 PORT MAP(
	A=> C(	1703	),
	B=>E(	1551	),
	Cin=> Carry( 	1638	),
	Cout=> Carry( 	1639	),
	S=> E(	1613	));
			
  U1640	: Somador_Exato_1 PORT MAP(
	A=> C(	1704	),
	B=>E(	1552	),
	Cin=> Carry( 	1639	),
	Cout=> Carry( 	1640	),
	S=> E(	1614	));
			
  U1641	: Somador_Exato_1 PORT MAP(
	A=> C(	1705	),
	B=>E(	1553	),
	Cin=> Carry( 	1640	),
	Cout=> Carry( 	1641	),
	S=> E(	1615	));
			
  U1642	: Somador_Exato_1 PORT MAP(
	A=> C(	1706	),
	B=>E(	1554	),
	Cin=> Carry( 	1641	),
	Cout=> Carry( 	1642	),
	S=> E(	1616	));
			
  U1643	: Somador_Exato_1 PORT MAP(
	A=> C(	1707	),
	B=>E(	1555	),
	Cin=> Carry( 	1642	),
	Cout=> Carry( 	1643	),
	S=> E(	1617	));
			
  U1644	: Somador_Exato_1 PORT MAP(
	A=> C(	1708	),
	B=>E(	1556	),
	Cin=> Carry( 	1643	),
	Cout=> Carry( 	1644	),
	S=> E(	1618	));
			
  U1645	: Somador_Exato_1 PORT MAP(
	A=> C(	1709	),
	B=>E(	1557	),
	Cin=> Carry( 	1644	),
	Cout=> Carry( 	1645	),
	S=> E(	1619	));
			
  U1646	: Somador_Exato_1 PORT MAP(
	A=> C(	1710	),
	B=>E(	1558	),
	Cin=> Carry( 	1645	),
	Cout=> Carry( 	1646	),
	S=> E(	1620	));
			
  U1647	: Somador_Exato_1 PORT MAP(
	A=> C(	1711	),
	B=>E(	1559	),
	Cin=> Carry( 	1646	),
	Cout=> Carry( 	1647	),
	S=> E(	1621	));
			
  U1648	: Somador_Exato_1 PORT MAP(
	A=> C(	1712	),
	B=>E(	1560	),
	Cin=> Carry( 	1647	),
	Cout=> Carry( 	1648	),
	S=> E(	1622	));
			
  U1649	: Somador_Exato_1 PORT MAP(
	A=> C(	1713	),
	B=>E(	1561	),
	Cin=> Carry( 	1648	),
	Cout=> Carry( 	1649	),
	S=> E(	1623	));
			
  U1650	: Somador_Exato_1 PORT MAP(
	A=> C(	1714	),
	B=>E(	1562	),
	Cin=> Carry( 	1649	),
	Cout=> Carry( 	1650	),
	S=> E(	1624	));
			
  U1651	: Somador_Exato_1 PORT MAP(
	A=> C(	1715	),
	B=>E(	1563	),
	Cin=> Carry( 	1650	),
	Cout=> Carry( 	1651	),
	S=> E(	1625	));
			
  U1652	: Somador_Exato_1 PORT MAP(
	A=> C(	1716	),
	B=>E(	1564	),
	Cin=> Carry( 	1651	),
	Cout=> Carry( 	1652	),
	S=> E(	1626	));
			
  U1653	: Somador_Exato_1 PORT MAP(
	A=> C(	1717	),
	B=>E(	1565	),
	Cin=> Carry( 	1652	),
	Cout=> Carry( 	1653	),
	S=> E(	1627	));
			
  U1654	: Somador_Exato_1 PORT MAP(
	A=> C(	1718	),
	B=>E(	1566	),
	Cin=> Carry( 	1653	),
	Cout=> Carry( 	1654	),
	S=> E(	1628	));
			
  U1655	: Somador_Exato_1 PORT MAP(
	A=> C(	1719	),
	B=>E(	1567	),
	Cin=> Carry( 	1654	),
	Cout=> Carry( 	1655	),
	S=> E(	1629	));
			
  U1656	: Somador_Exato_1 PORT MAP(
	A=> C(	1720	),
	B=>E(	1568	),
	Cin=> Carry( 	1655	),
	Cout=> Carry( 	1656	),
	S=> E(	1630	));
			
  U1657	: Somador_Exato_1 PORT MAP(
	A=> C(	1721	),
	B=>E(	1569	),
	Cin=> Carry( 	1656	),
	Cout=> Carry( 	1657	),
	S=> E(	1631	));
			
  U1658	: Somador_Exato_1 PORT MAP(
	A=> C(	1722	),
	B=>E(	1570	),
	Cin=> Carry( 	1657	),
	Cout=> Carry( 	1658	),
	S=> E(	1632	));
			
  U1659	: Somador_Exato_1 PORT MAP(
	A=> C(	1723	),
	B=>E(	1571	),
	Cin=> Carry( 	1658	),
	Cout=> Carry( 	1659	),
	S=> E(	1633	));
			
  U1660	: Somador_Exato_1 PORT MAP(
	A=> C(	1724	),
	B=>E(	1572	),
	Cin=> Carry( 	1659	),
	Cout=> Carry( 	1660	),
	S=> E(	1634	));
			
  U1661	: Somador_Exato_1 PORT MAP(
	A=> C(	1725	),
	B=>E(	1573	),
	Cin=> Carry( 	1660	),
	Cout=> Carry( 	1661	),
	S=> E(	1635	));
			
  U1662	: Somador_Exato_1 PORT MAP(
	A=> C(	1726	),
	B=>E(	1574	),
	Cin=> Carry( 	1661	),
	Cout=> Carry( 	1662	),
	S=> E(	1636	));
			
  U1663	: Somador_Exato_1 PORT MAP(
	A=> C(	1727	),
	B=>Carry(	1599	),
	Cin=> Carry( 	1662	),
	Cout=> Carry( 	1663	),
	S=> E(	1637	));

			
  U1664	: Somador_Exato_1 PORT MAP(
	A=> C(	1728	),
	B=>E(	1575	),
	Cin=> '0'	,
	Cout=> Carry( 	1664	),
	S=> R(	27	));
			
  U1665	: Somador_Exato_1 PORT MAP(
	A=> C(	1729	),
	B=>E(	1576	),
	Cin=> Carry( 	1664	),
	Cout=> Carry( 	1665	),
	S=> E(	1638	));
			
  U1666	: Somador_Exato_1 PORT MAP(
	A=> C(	1730	),
	B=>E(	1577	),
	Cin=> Carry( 	1665	),
	Cout=> Carry( 	1666	),
	S=> E(	1639	));
			
  U1667	: Somador_Exato_1 PORT MAP(
	A=> C(	1731	),
	B=>E(	1578	),
	Cin=> Carry( 	1666	),
	Cout=> Carry( 	1667	),
	S=> E(	1640	));
			
  U1668	: Somador_Exato_1 PORT MAP(
	A=> C(	1732	),
	B=>E(	1579	),
	Cin=> Carry( 	1667	),
	Cout=> Carry( 	1668	),
	S=> E(	1641	));
			
  U1669	: Somador_Exato_1 PORT MAP(
	A=> C(	1733	),
	B=>E(	1580	),
	Cin=> Carry( 	1668	),
	Cout=> Carry( 	1669	),
	S=> E(	1642	));
			
  U1670	: Somador_Exato_1 PORT MAP(
	A=> C(	1734	),
	B=>E(	1581	),
	Cin=> Carry( 	1669	),
	Cout=> Carry( 	1670	),
	S=> E(	1643	));
			
  U1671	: Somador_Exato_1 PORT MAP(
	A=> C(	1735	),
	B=>E(	1582	),
	Cin=> Carry( 	1670	),
	Cout=> Carry( 	1671	),
	S=> E(	1644	));
			
  U1672	: Somador_Exato_1 PORT MAP(
	A=> C(	1736	),
	B=>E(	1583	),
	Cin=> Carry( 	1671	),
	Cout=> Carry( 	1672	),
	S=> E(	1645	));
			
  U1673	: Somador_Exato_1 PORT MAP(
	A=> C(	1737	),
	B=>E(	1584	),
	Cin=> Carry( 	1672	),
	Cout=> Carry( 	1673	),
	S=> E(	1646	));
			
  U1674	: Somador_Exato_1 PORT MAP(
	A=> C(	1738	),
	B=>E(	1585	),
	Cin=> Carry( 	1673	),
	Cout=> Carry( 	1674	),
	S=> E(	1647	));
			
  U1675	: Somador_Exato_1 PORT MAP(
	A=> C(	1739	),
	B=>E(	1586	),
	Cin=> Carry( 	1674	),
	Cout=> Carry( 	1675	),
	S=> E(	1648	));
			
  U1676	: Somador_Exato_1 PORT MAP(
	A=> C(	1740	),
	B=>E(	1587	),
	Cin=> Carry( 	1675	),
	Cout=> Carry( 	1676	),
	S=> E(	1649	));
			
  U1677	: Somador_Exato_1 PORT MAP(
	A=> C(	1741	),
	B=>E(	1588	),
	Cin=> Carry( 	1676	),
	Cout=> Carry( 	1677	),
	S=> E(	1650	));
			
  U1678	: Somador_Exato_1 PORT MAP(
	A=> C(	1742	),
	B=>E(	1589	),
	Cin=> Carry( 	1677	),
	Cout=> Carry( 	1678	),
	S=> E(	1651	));
			
  U1679	: Somador_Exato_1 PORT MAP(
	A=> C(	1743	),
	B=>E(	1590	),
	Cin=> Carry( 	1678	),
	Cout=> Carry( 	1679	),
	S=> E(	1652	));
			
  U1680	: Somador_Exato_1 PORT MAP(
	A=> C(	1744	),
	B=>E(	1591	),
	Cin=> Carry( 	1679	),
	Cout=> Carry( 	1680	),
	S=> E(	1653	));
			
  U1681	: Somador_Exato_1 PORT MAP(
	A=> C(	1745	),
	B=>E(	1592	),
	Cin=> Carry( 	1680	),
	Cout=> Carry( 	1681	),
	S=> E(	1654	));
			
  U1682	: Somador_Exato_1 PORT MAP(
	A=> C(	1746	),
	B=>E(	1593	),
	Cin=> Carry( 	1681	),
	Cout=> Carry( 	1682	),
	S=> E(	1655	));
			
  U1683	: Somador_Exato_1 PORT MAP(
	A=> C(	1747	),
	B=>E(	1594	),
	Cin=> Carry( 	1682	),
	Cout=> Carry( 	1683	),
	S=> E(	1656	));
			
  U1684	: Somador_Exato_1 PORT MAP(
	A=> C(	1748	),
	B=>E(	1595	),
	Cin=> Carry( 	1683	),
	Cout=> Carry( 	1684	),
	S=> E(	1657	));
			
  U1685	: Somador_Exato_1 PORT MAP(
	A=> C(	1749	),
	B=>E(	1596	),
	Cin=> Carry( 	1684	),
	Cout=> Carry( 	1685	),
	S=> E(	1658	));
			
  U1686	: Somador_Exato_1 PORT MAP(
	A=> C(	1750	),
	B=>E(	1597	),
	Cin=> Carry( 	1685	),
	Cout=> Carry( 	1686	),
	S=> E(	1659	));
			
  U1687	: Somador_Exato_1 PORT MAP(
	A=> C(	1751	),
	B=>E(	1598	),
	Cin=> Carry( 	1686	),
	Cout=> Carry( 	1687	),
	S=> E(	1660	));
			
  U1688	: Somador_Exato_1 PORT MAP(
	A=> C(	1752	),
	B=>E(	1599	),
	Cin=> Carry( 	1687	),
	Cout=> Carry( 	1688	),
	S=> E(	1661	));
			
  U1689	: Somador_Exato_1 PORT MAP(
	A=> C(	1753	),
	B=>E(	1600	),
	Cin=> Carry( 	1688	),
	Cout=> Carry( 	1689	),
	S=> E(	1662	));
			
  U1690	: Somador_Exato_1 PORT MAP(
	A=> C(	1754	),
	B=>E(	1601	),
	Cin=> Carry( 	1689	),
	Cout=> Carry( 	1690	),
	S=> E(	1663	));
			
  U1691	: Somador_Exato_1 PORT MAP(
	A=> C(	1755	),
	B=>E(	1602	),
	Cin=> Carry( 	1690	),
	Cout=> Carry( 	1691	),
	S=> E(	1664	));
			
  U1692	: Somador_Exato_1 PORT MAP(
	A=> C(	1756	),
	B=>E(	1603	),
	Cin=> Carry( 	1691	),
	Cout=> Carry( 	1692	),
	S=> E(	1665	));
			
  U1693	: Somador_Exato_1 PORT MAP(
	A=> C(	1757	),
	B=>E(	1604	),
	Cin=> Carry( 	1692	),
	Cout=> Carry( 	1693	),
	S=> E(	1666	));
			
  U1694	: Somador_Exato_1 PORT MAP(
	A=> C(	1758	),
	B=>E(	1605	),
	Cin=> Carry( 	1693	),
	Cout=> Carry( 	1694	),
	S=> E(	1667	));
			
  U1695	: Somador_Exato_1 PORT MAP(
	A=> C(	1759	),
	B=>E(	1606	),
	Cin=> Carry( 	1694	),
	Cout=> Carry( 	1695	),
	S=> E(	1668	));
			
  U1696	: Somador_Exato_1 PORT MAP(
	A=> C(	1760	),
	B=>E(	1607	),
	Cin=> Carry( 	1695	),
	Cout=> Carry( 	1696	),
	S=> E(	1669	));
			
  U1697	: Somador_Exato_1 PORT MAP(
	A=> C(	1761	),
	B=>E(	1608	),
	Cin=> Carry( 	1696	),
	Cout=> Carry( 	1697	),
	S=> E(	1670	));
			
  U1698	: Somador_Exato_1 PORT MAP(
	A=> C(	1762	),
	B=>E(	1609	),
	Cin=> Carry( 	1697	),
	Cout=> Carry( 	1698	),
	S=> E(	1671	));
			
  U1699	: Somador_Exato_1 PORT MAP(
	A=> C(	1763	),
	B=>E(	1610	),
	Cin=> Carry( 	1698	),
	Cout=> Carry( 	1699	),
	S=> E(	1672	));
			
  U1700	: Somador_Exato_1 PORT MAP(
	A=> C(	1764	),
	B=>E(	1611	),
	Cin=> Carry( 	1699	),
	Cout=> Carry( 	1700	),
	S=> E(	1673	));
			
  U1701	: Somador_Exato_1 PORT MAP(
	A=> C(	1765	),
	B=>E(	1612	),
	Cin=> Carry( 	1700	),
	Cout=> Carry( 	1701	),
	S=> E(	1674	));
			
  U1702	: Somador_Exato_1 PORT MAP(
	A=> C(	1766	),
	B=>E(	1613	),
	Cin=> Carry( 	1701	),
	Cout=> Carry( 	1702	),
	S=> E(	1675	));
			
  U1703	: Somador_Exato_1 PORT MAP(
	A=> C(	1767	),
	B=>E(	1614	),
	Cin=> Carry( 	1702	),
	Cout=> Carry( 	1703	),
	S=> E(	1676	));
			
  U1704	: Somador_Exato_1 PORT MAP(
	A=> C(	1768	),
	B=>E(	1615	),
	Cin=> Carry( 	1703	),
	Cout=> Carry( 	1704	),
	S=> E(	1677	));
			
  U1705	: Somador_Exato_1 PORT MAP(
	A=> C(	1769	),
	B=>E(	1616	),
	Cin=> Carry( 	1704	),
	Cout=> Carry( 	1705	),
	S=> E(	1678	));
			
  U1706	: Somador_Exato_1 PORT MAP(
	A=> C(	1770	),
	B=>E(	1617	),
	Cin=> Carry( 	1705	),
	Cout=> Carry( 	1706	),
	S=> E(	1679	));
			
  U1707	: Somador_Exato_1 PORT MAP(
	A=> C(	1771	),
	B=>E(	1618	),
	Cin=> Carry( 	1706	),
	Cout=> Carry( 	1707	),
	S=> E(	1680	));
			
  U1708	: Somador_Exato_1 PORT MAP(
	A=> C(	1772	),
	B=>E(	1619	),
	Cin=> Carry( 	1707	),
	Cout=> Carry( 	1708	),
	S=> E(	1681	));
			
  U1709	: Somador_Exato_1 PORT MAP(
	A=> C(	1773	),
	B=>E(	1620	),
	Cin=> Carry( 	1708	),
	Cout=> Carry( 	1709	),
	S=> E(	1682	));
			
  U1710	: Somador_Exato_1 PORT MAP(
	A=> C(	1774	),
	B=>E(	1621	),
	Cin=> Carry( 	1709	),
	Cout=> Carry( 	1710	),
	S=> E(	1683	));
			
  U1711	: Somador_Exato_1 PORT MAP(
	A=> C(	1775	),
	B=>E(	1622	),
	Cin=> Carry( 	1710	),
	Cout=> Carry( 	1711	),
	S=> E(	1684	));
			
  U1712	: Somador_Exato_1 PORT MAP(
	A=> C(	1776	),
	B=>E(	1623	),
	Cin=> Carry( 	1711	),
	Cout=> Carry( 	1712	),
	S=> E(	1685	));
			
  U1713	: Somador_Exato_1 PORT MAP(
	A=> C(	1777	),
	B=>E(	1624	),
	Cin=> Carry( 	1712	),
	Cout=> Carry( 	1713	),
	S=> E(	1686	));
			
  U1714	: Somador_Exato_1 PORT MAP(
	A=> C(	1778	),
	B=>E(	1625	),
	Cin=> Carry( 	1713	),
	Cout=> Carry( 	1714	),
	S=> E(	1687	));
			
  U1715	: Somador_Exato_1 PORT MAP(
	A=> C(	1779	),
	B=>E(	1626	),
	Cin=> Carry( 	1714	),
	Cout=> Carry( 	1715	),
	S=> E(	1688	));
			
  U1716	: Somador_Exato_1 PORT MAP(
	A=> C(	1780	),
	B=>E(	1627	),
	Cin=> Carry( 	1715	),
	Cout=> Carry( 	1716	),
	S=> E(	1689	));
			
  U1717	: Somador_Exato_1 PORT MAP(
	A=> C(	1781	),
	B=>E(	1628	),
	Cin=> Carry( 	1716	),
	Cout=> Carry( 	1717	),
	S=> E(	1690	));
			
  U1718	: Somador_Exato_1 PORT MAP(
	A=> C(	1782	),
	B=>E(	1629	),
	Cin=> Carry( 	1717	),
	Cout=> Carry( 	1718	),
	S=> E(	1691	));
			
  U1719	: Somador_Exato_1 PORT MAP(
	A=> C(	1783	),
	B=>E(	1630	),
	Cin=> Carry( 	1718	),
	Cout=> Carry( 	1719	),
	S=> E(	1692	));
			
  U1720	: Somador_Exato_1 PORT MAP(
	A=> C(	1784	),
	B=>E(	1631	),
	Cin=> Carry( 	1719	),
	Cout=> Carry( 	1720	),
	S=> E(	1693	));
			
  U1721	: Somador_Exato_1 PORT MAP(
	A=> C(	1785	),
	B=>E(	1632	),
	Cin=> Carry( 	1720	),
	Cout=> Carry( 	1721	),
	S=> E(	1694	));
			
  U1722	: Somador_Exato_1 PORT MAP(
	A=> C(	1786	),
	B=>E(	1633	),
	Cin=> Carry( 	1721	),
	Cout=> Carry( 	1722	),
	S=> E(	1695	));
			
  U1723	: Somador_Exato_1 PORT MAP(
	A=> C(	1787	),
	B=>E(	1634	),
	Cin=> Carry( 	1722	),
	Cout=> Carry( 	1723	),
	S=> E(	1696	));
			
  U1724	: Somador_Exato_1 PORT MAP(
	A=> C(	1788	),
	B=>E(	1635	),
	Cin=> Carry( 	1723	),
	Cout=> Carry( 	1724	),
	S=> E(	1697	));
			
  U1725	: Somador_Exato_1 PORT MAP(
	A=> C(	1789	),
	B=>E(	1636	),
	Cin=> Carry( 	1724	),
	Cout=> Carry( 	1725	),
	S=> E(	1698	));
			
  U1726	: Somador_Exato_1 PORT MAP(
	A=> C(	1790	),
	B=>E(	1637	),
	Cin=> Carry( 	1725	),
	Cout=> Carry( 	1726	),
	S=> E(	1699	));
			
  U1727	: Somador_Exato_1 PORT MAP(
	A=> C(	1791	),
	B=>Carry(	1663	),
	Cin=> Carry( 	1726	),
	Cout=> Carry( 	1727	),
	S=> E(	1700	));

			
  U1728	: Somador_Exato_1 PORT MAP(
	A=> C(	1792	),
	B=>E(	1638	),
	Cin=> '0'	,
	Cout=> Carry( 	1728	),
	S=> R(	28	));
			
  U1729	: Somador_Exato_1 PORT MAP(
	A=> C(	1793	),
	B=>E(	1639	),
	Cin=> Carry( 	1728	),
	Cout=> Carry( 	1729	),
	S=> E(	1701	));
			
  U1730	: Somador_Exato_1 PORT MAP(
	A=> C(	1794	),
	B=>E(	1640	),
	Cin=> Carry( 	1729	),
	Cout=> Carry( 	1730	),
	S=> E(	1702	));
			
  U1731	: Somador_Exato_1 PORT MAP(
	A=> C(	1795	),
	B=>E(	1641	),
	Cin=> Carry( 	1730	),
	Cout=> Carry( 	1731	),
	S=> E(	1703	));
			
  U1732	: Somador_Exato_1 PORT MAP(
	A=> C(	1796	),
	B=>E(	1642	),
	Cin=> Carry( 	1731	),
	Cout=> Carry( 	1732	),
	S=> E(	1704	));
			
  U1733	: Somador_Exato_1 PORT MAP(
	A=> C(	1797	),
	B=>E(	1643	),
	Cin=> Carry( 	1732	),
	Cout=> Carry( 	1733	),
	S=> E(	1705	));
			
  U1734	: Somador_Exato_1 PORT MAP(
	A=> C(	1798	),
	B=>E(	1644	),
	Cin=> Carry( 	1733	),
	Cout=> Carry( 	1734	),
	S=> E(	1706	));
			
  U1735	: Somador_Exato_1 PORT MAP(
	A=> C(	1799	),
	B=>E(	1645	),
	Cin=> Carry( 	1734	),
	Cout=> Carry( 	1735	),
	S=> E(	1707	));
			
  U1736	: Somador_Exato_1 PORT MAP(
	A=> C(	1800	),
	B=>E(	1646	),
	Cin=> Carry( 	1735	),
	Cout=> Carry( 	1736	),
	S=> E(	1708	));
			
  U1737	: Somador_Exato_1 PORT MAP(
	A=> C(	1801	),
	B=>E(	1647	),
	Cin=> Carry( 	1736	),
	Cout=> Carry( 	1737	),
	S=> E(	1709	));
			
  U1738	: Somador_Exato_1 PORT MAP(
	A=> C(	1802	),
	B=>E(	1648	),
	Cin=> Carry( 	1737	),
	Cout=> Carry( 	1738	),
	S=> E(	1710	));
			
  U1739	: Somador_Exato_1 PORT MAP(
	A=> C(	1803	),
	B=>E(	1649	),
	Cin=> Carry( 	1738	),
	Cout=> Carry( 	1739	),
	S=> E(	1711	));
			
  U1740	: Somador_Exato_1 PORT MAP(
	A=> C(	1804	),
	B=>E(	1650	),
	Cin=> Carry( 	1739	),
	Cout=> Carry( 	1740	),
	S=> E(	1712	));
			
  U1741	: Somador_Exato_1 PORT MAP(
	A=> C(	1805	),
	B=>E(	1651	),
	Cin=> Carry( 	1740	),
	Cout=> Carry( 	1741	),
	S=> E(	1713	));
			
  U1742	: Somador_Exato_1 PORT MAP(
	A=> C(	1806	),
	B=>E(	1652	),
	Cin=> Carry( 	1741	),
	Cout=> Carry( 	1742	),
	S=> E(	1714	));
			
  U1743	: Somador_Exato_1 PORT MAP(
	A=> C(	1807	),
	B=>E(	1653	),
	Cin=> Carry( 	1742	),
	Cout=> Carry( 	1743	),
	S=> E(	1715	));
			
  U1744	: Somador_Exato_1 PORT MAP(
	A=> C(	1808	),
	B=>E(	1654	),
	Cin=> Carry( 	1743	),
	Cout=> Carry( 	1744	),
	S=> E(	1716	));
			
  U1745	: Somador_Exato_1 PORT MAP(
	A=> C(	1809	),
	B=>E(	1655	),
	Cin=> Carry( 	1744	),
	Cout=> Carry( 	1745	),
	S=> E(	1717	));
			
  U1746	: Somador_Exato_1 PORT MAP(
	A=> C(	1810	),
	B=>E(	1656	),
	Cin=> Carry( 	1745	),
	Cout=> Carry( 	1746	),
	S=> E(	1718	));
			
  U1747	: Somador_Exato_1 PORT MAP(
	A=> C(	1811	),
	B=>E(	1657	),
	Cin=> Carry( 	1746	),
	Cout=> Carry( 	1747	),
	S=> E(	1719	));
			
  U1748	: Somador_Exato_1 PORT MAP(
	A=> C(	1812	),
	B=>E(	1658	),
	Cin=> Carry( 	1747	),
	Cout=> Carry( 	1748	),
	S=> E(	1720	));
			
  U1749	: Somador_Exato_1 PORT MAP(
	A=> C(	1813	),
	B=>E(	1659	),
	Cin=> Carry( 	1748	),
	Cout=> Carry( 	1749	),
	S=> E(	1721	));
			
  U1750	: Somador_Exato_1 PORT MAP(
	A=> C(	1814	),
	B=>E(	1660	),
	Cin=> Carry( 	1749	),
	Cout=> Carry( 	1750	),
	S=> E(	1722	));
			
  U1751	: Somador_Exato_1 PORT MAP(
	A=> C(	1815	),
	B=>E(	1661	),
	Cin=> Carry( 	1750	),
	Cout=> Carry( 	1751	),
	S=> E(	1723	));
			
  U1752	: Somador_Exato_1 PORT MAP(
	A=> C(	1816	),
	B=>E(	1662	),
	Cin=> Carry( 	1751	),
	Cout=> Carry( 	1752	),
	S=> E(	1724	));
			
  U1753	: Somador_Exato_1 PORT MAP(
	A=> C(	1817	),
	B=>E(	1663	),
	Cin=> Carry( 	1752	),
	Cout=> Carry( 	1753	),
	S=> E(	1725	));
			
  U1754	: Somador_Exato_1 PORT MAP(
	A=> C(	1818	),
	B=>E(	1664	),
	Cin=> Carry( 	1753	),
	Cout=> Carry( 	1754	),
	S=> E(	1726	));
			
  U1755	: Somador_Exato_1 PORT MAP(
	A=> C(	1819	),
	B=>E(	1665	),
	Cin=> Carry( 	1754	),
	Cout=> Carry( 	1755	),
	S=> E(	1727	));
			
  U1756	: Somador_Exato_1 PORT MAP(
	A=> C(	1820	),
	B=>E(	1666	),
	Cin=> Carry( 	1755	),
	Cout=> Carry( 	1756	),
	S=> E(	1728	));
			
  U1757	: Somador_Exato_1 PORT MAP(
	A=> C(	1821	),
	B=>E(	1667	),
	Cin=> Carry( 	1756	),
	Cout=> Carry( 	1757	),
	S=> E(	1729	));
			
  U1758	: Somador_Exato_1 PORT MAP(
	A=> C(	1822	),
	B=>E(	1668	),
	Cin=> Carry( 	1757	),
	Cout=> Carry( 	1758	),
	S=> E(	1730	));
			
  U1759	: Somador_Exato_1 PORT MAP(
	A=> C(	1823	),
	B=>E(	1669	),
	Cin=> Carry( 	1758	),
	Cout=> Carry( 	1759	),
	S=> E(	1731	));
			
  U1760	: Somador_Exato_1 PORT MAP(
	A=> C(	1824	),
	B=>E(	1670	),
	Cin=> Carry( 	1759	),
	Cout=> Carry( 	1760	),
	S=> E(	1732	));
			
  U1761	: Somador_Exato_1 PORT MAP(
	A=> C(	1825	),
	B=>E(	1671	),
	Cin=> Carry( 	1760	),
	Cout=> Carry( 	1761	),
	S=> E(	1733	));
			
  U1762	: Somador_Exato_1 PORT MAP(
	A=> C(	1826	),
	B=>E(	1672	),
	Cin=> Carry( 	1761	),
	Cout=> Carry( 	1762	),
	S=> E(	1734	));
			
  U1763	: Somador_Exato_1 PORT MAP(
	A=> C(	1827	),
	B=>E(	1673	),
	Cin=> Carry( 	1762	),
	Cout=> Carry( 	1763	),
	S=> E(	1735	));
			
  U1764	: Somador_Exato_1 PORT MAP(
	A=> C(	1828	),
	B=>E(	1674	),
	Cin=> Carry( 	1763	),
	Cout=> Carry( 	1764	),
	S=> E(	1736	));
			
  U1765	: Somador_Exato_1 PORT MAP(
	A=> C(	1829	),
	B=>E(	1675	),
	Cin=> Carry( 	1764	),
	Cout=> Carry( 	1765	),
	S=> E(	1737	));
			
  U1766	: Somador_Exato_1 PORT MAP(
	A=> C(	1830	),
	B=>E(	1676	),
	Cin=> Carry( 	1765	),
	Cout=> Carry( 	1766	),
	S=> E(	1738	));
			
  U1767	: Somador_Exato_1 PORT MAP(
	A=> C(	1831	),
	B=>E(	1677	),
	Cin=> Carry( 	1766	),
	Cout=> Carry( 	1767	),
	S=> E(	1739	));
			
  U1768	: Somador_Exato_1 PORT MAP(
	A=> C(	1832	),
	B=>E(	1678	),
	Cin=> Carry( 	1767	),
	Cout=> Carry( 	1768	),
	S=> E(	1740	));
			
  U1769	: Somador_Exato_1 PORT MAP(
	A=> C(	1833	),
	B=>E(	1679	),
	Cin=> Carry( 	1768	),
	Cout=> Carry( 	1769	),
	S=> E(	1741	));
			
  U1770	: Somador_Exato_1 PORT MAP(
	A=> C(	1834	),
	B=>E(	1680	),
	Cin=> Carry( 	1769	),
	Cout=> Carry( 	1770	),
	S=> E(	1742	));
			
  U1771	: Somador_Exato_1 PORT MAP(
	A=> C(	1835	),
	B=>E(	1681	),
	Cin=> Carry( 	1770	),
	Cout=> Carry( 	1771	),
	S=> E(	1743	));
			
  U1772	: Somador_Exato_1 PORT MAP(
	A=> C(	1836	),
	B=>E(	1682	),
	Cin=> Carry( 	1771	),
	Cout=> Carry( 	1772	),
	S=> E(	1744	));
			
  U1773	: Somador_Exato_1 PORT MAP(
	A=> C(	1837	),
	B=>E(	1683	),
	Cin=> Carry( 	1772	),
	Cout=> Carry( 	1773	),
	S=> E(	1745	));
			
  U1774	: Somador_Exato_1 PORT MAP(
	A=> C(	1838	),
	B=>E(	1684	),
	Cin=> Carry( 	1773	),
	Cout=> Carry( 	1774	),
	S=> E(	1746	));
			
  U1775	: Somador_Exato_1 PORT MAP(
	A=> C(	1839	),
	B=>E(	1685	),
	Cin=> Carry( 	1774	),
	Cout=> Carry( 	1775	),
	S=> E(	1747	));
			
  U1776	: Somador_Exato_1 PORT MAP(
	A=> C(	1840	),
	B=>E(	1686	),
	Cin=> Carry( 	1775	),
	Cout=> Carry( 	1776	),
	S=> E(	1748	));
			
  U1777	: Somador_Exato_1 PORT MAP(
	A=> C(	1841	),
	B=>E(	1687	),
	Cin=> Carry( 	1776	),
	Cout=> Carry( 	1777	),
	S=> E(	1749	));
			
  U1778	: Somador_Exato_1 PORT MAP(
	A=> C(	1842	),
	B=>E(	1688	),
	Cin=> Carry( 	1777	),
	Cout=> Carry( 	1778	),
	S=> E(	1750	));
			
  U1779	: Somador_Exato_1 PORT MAP(
	A=> C(	1843	),
	B=>E(	1689	),
	Cin=> Carry( 	1778	),
	Cout=> Carry( 	1779	),
	S=> E(	1751	));
			
  U1780	: Somador_Exato_1 PORT MAP(
	A=> C(	1844	),
	B=>E(	1690	),
	Cin=> Carry( 	1779	),
	Cout=> Carry( 	1780	),
	S=> E(	1752	));
			
  U1781	: Somador_Exato_1 PORT MAP(
	A=> C(	1845	),
	B=>E(	1691	),
	Cin=> Carry( 	1780	),
	Cout=> Carry( 	1781	),
	S=> E(	1753	));
			
  U1782	: Somador_Exato_1 PORT MAP(
	A=> C(	1846	),
	B=>E(	1692	),
	Cin=> Carry( 	1781	),
	Cout=> Carry( 	1782	),
	S=> E(	1754	));
			
  U1783	: Somador_Exato_1 PORT MAP(
	A=> C(	1847	),
	B=>E(	1693	),
	Cin=> Carry( 	1782	),
	Cout=> Carry( 	1783	),
	S=> E(	1755	));
			
  U1784	: Somador_Exato_1 PORT MAP(
	A=> C(	1848	),
	B=>E(	1694	),
	Cin=> Carry( 	1783	),
	Cout=> Carry( 	1784	),
	S=> E(	1756	));
			
  U1785	: Somador_Exato_1 PORT MAP(
	A=> C(	1849	),
	B=>E(	1695	),
	Cin=> Carry( 	1784	),
	Cout=> Carry( 	1785	),
	S=> E(	1757	));
			
  U1786	: Somador_Exato_1 PORT MAP(
	A=> C(	1850	),
	B=>E(	1696	),
	Cin=> Carry( 	1785	),
	Cout=> Carry( 	1786	),
	S=> E(	1758	));
			
  U1787	: Somador_Exato_1 PORT MAP(
	A=> C(	1851	),
	B=>E(	1697	),
	Cin=> Carry( 	1786	),
	Cout=> Carry( 	1787	),
	S=> E(	1759	));
			
  U1788	: Somador_Exato_1 PORT MAP(
	A=> C(	1852	),
	B=>E(	1698	),
	Cin=> Carry( 	1787	),
	Cout=> Carry( 	1788	),
	S=> E(	1760	));
			
  U1789	: Somador_Exato_1 PORT MAP(
	A=> C(	1853	),
	B=>E(	1699	),
	Cin=> Carry( 	1788	),
	Cout=> Carry( 	1789	),
	S=> E(	1761	));
			
  U1790	: Somador_Exato_1 PORT MAP(
	A=> C(	1854	),
	B=>E(	1700	),
	Cin=> Carry( 	1789	),
	Cout=> Carry( 	1790	),
	S=> E(	1762	));
			
  U1791	: Somador_Exato_1 PORT MAP(
	A=> C(	1855	),
	B=>Carry(	1727	),
	Cin=> Carry( 	1790	),
	Cout=> Carry( 	1791	),
	S=> E(	1763	));

			
  U1792	: Somador_Exato_1 PORT MAP(
	A=> C(	1856	),
	B=>E(	1701	),
	Cin=> '0'	,
	Cout=> Carry( 	1792	),
	S=> R(	29	));
			
  U1793	: Somador_Exato_1 PORT MAP(
	A=> C(	1857	),
	B=>E(	1702	),
	Cin=> Carry( 	1792	),
	Cout=> Carry( 	1793	),
	S=> E(	1764	));
			
  U1794	: Somador_Exato_1 PORT MAP(
	A=> C(	1858	),
	B=>E(	1703	),
	Cin=> Carry( 	1793	),
	Cout=> Carry( 	1794	),
	S=> E(	1765	));
			
  U1795	: Somador_Exato_1 PORT MAP(
	A=> C(	1859	),
	B=>E(	1704	),
	Cin=> Carry( 	1794	),
	Cout=> Carry( 	1795	),
	S=> E(	1766	));
			
  U1796	: Somador_Exato_1 PORT MAP(
	A=> C(	1860	),
	B=>E(	1705	),
	Cin=> Carry( 	1795	),
	Cout=> Carry( 	1796	),
	S=> E(	1767	));
			
  U1797	: Somador_Exato_1 PORT MAP(
	A=> C(	1861	),
	B=>E(	1706	),
	Cin=> Carry( 	1796	),
	Cout=> Carry( 	1797	),
	S=> E(	1768	));
			
  U1798	: Somador_Exato_1 PORT MAP(
	A=> C(	1862	),
	B=>E(	1707	),
	Cin=> Carry( 	1797	),
	Cout=> Carry( 	1798	),
	S=> E(	1769	));
			
  U1799	: Somador_Exato_1 PORT MAP(
	A=> C(	1863	),
	B=>E(	1708	),
	Cin=> Carry( 	1798	),
	Cout=> Carry( 	1799	),
	S=> E(	1770	));
			
  U1800	: Somador_Exato_1 PORT MAP(
	A=> C(	1864	),
	B=>E(	1709	),
	Cin=> Carry( 	1799	),
	Cout=> Carry( 	1800	),
	S=> E(	1771	));
			
  U1801	: Somador_Exato_1 PORT MAP(
	A=> C(	1865	),
	B=>E(	1710	),
	Cin=> Carry( 	1800	),
	Cout=> Carry( 	1801	),
	S=> E(	1772	));
			
  U1802	: Somador_Exato_1 PORT MAP(
	A=> C(	1866	),
	B=>E(	1711	),
	Cin=> Carry( 	1801	),
	Cout=> Carry( 	1802	),
	S=> E(	1773	));
			
  U1803	: Somador_Exato_1 PORT MAP(
	A=> C(	1867	),
	B=>E(	1712	),
	Cin=> Carry( 	1802	),
	Cout=> Carry( 	1803	),
	S=> E(	1774	));
			
  U1804	: Somador_Exato_1 PORT MAP(
	A=> C(	1868	),
	B=>E(	1713	),
	Cin=> Carry( 	1803	),
	Cout=> Carry( 	1804	),
	S=> E(	1775	));
			
  U1805	: Somador_Exato_1 PORT MAP(
	A=> C(	1869	),
	B=>E(	1714	),
	Cin=> Carry( 	1804	),
	Cout=> Carry( 	1805	),
	S=> E(	1776	));
			
  U1806	: Somador_Exato_1 PORT MAP(
	A=> C(	1870	),
	B=>E(	1715	),
	Cin=> Carry( 	1805	),
	Cout=> Carry( 	1806	),
	S=> E(	1777	));
			
  U1807	: Somador_Exato_1 PORT MAP(
	A=> C(	1871	),
	B=>E(	1716	),
	Cin=> Carry( 	1806	),
	Cout=> Carry( 	1807	),
	S=> E(	1778	));
			
  U1808	: Somador_Exato_1 PORT MAP(
	A=> C(	1872	),
	B=>E(	1717	),
	Cin=> Carry( 	1807	),
	Cout=> Carry( 	1808	),
	S=> E(	1779	));
			
  U1809	: Somador_Exato_1 PORT MAP(
	A=> C(	1873	),
	B=>E(	1718	),
	Cin=> Carry( 	1808	),
	Cout=> Carry( 	1809	),
	S=> E(	1780	));
			
  U1810	: Somador_Exato_1 PORT MAP(
	A=> C(	1874	),
	B=>E(	1719	),
	Cin=> Carry( 	1809	),
	Cout=> Carry( 	1810	),
	S=> E(	1781	));
			
  U1811	: Somador_Exato_1 PORT MAP(
	A=> C(	1875	),
	B=>E(	1720	),
	Cin=> Carry( 	1810	),
	Cout=> Carry( 	1811	),
	S=> E(	1782	));
			
  U1812	: Somador_Exato_1 PORT MAP(
	A=> C(	1876	),
	B=>E(	1721	),
	Cin=> Carry( 	1811	),
	Cout=> Carry( 	1812	),
	S=> E(	1783	));
			
  U1813	: Somador_Exato_1 PORT MAP(
	A=> C(	1877	),
	B=>E(	1722	),
	Cin=> Carry( 	1812	),
	Cout=> Carry( 	1813	),
	S=> E(	1784	));
			
  U1814	: Somador_Exato_1 PORT MAP(
	A=> C(	1878	),
	B=>E(	1723	),
	Cin=> Carry( 	1813	),
	Cout=> Carry( 	1814	),
	S=> E(	1785	));
			
  U1815	: Somador_Exato_1 PORT MAP(
	A=> C(	1879	),
	B=>E(	1724	),
	Cin=> Carry( 	1814	),
	Cout=> Carry( 	1815	),
	S=> E(	1786	));
			
  U1816	: Somador_Exato_1 PORT MAP(
	A=> C(	1880	),
	B=>E(	1725	),
	Cin=> Carry( 	1815	),
	Cout=> Carry( 	1816	),
	S=> E(	1787	));
			
  U1817	: Somador_Exato_1 PORT MAP(
	A=> C(	1881	),
	B=>E(	1726	),
	Cin=> Carry( 	1816	),
	Cout=> Carry( 	1817	),
	S=> E(	1788	));
			
  U1818	: Somador_Exato_1 PORT MAP(
	A=> C(	1882	),
	B=>E(	1727	),
	Cin=> Carry( 	1817	),
	Cout=> Carry( 	1818	),
	S=> E(	1789	));
			
  U1819	: Somador_Exato_1 PORT MAP(
	A=> C(	1883	),
	B=>E(	1728	),
	Cin=> Carry( 	1818	),
	Cout=> Carry( 	1819	),
	S=> E(	1790	));
			
  U1820	: Somador_Exato_1 PORT MAP(
	A=> C(	1884	),
	B=>E(	1729	),
	Cin=> Carry( 	1819	),
	Cout=> Carry( 	1820	),
	S=> E(	1791	));
			
  U1821	: Somador_Exato_1 PORT MAP(
	A=> C(	1885	),
	B=>E(	1730	),
	Cin=> Carry( 	1820	),
	Cout=> Carry( 	1821	),
	S=> E(	1792	));
			
  U1822	: Somador_Exato_1 PORT MAP(
	A=> C(	1886	),
	B=>E(	1731	),
	Cin=> Carry( 	1821	),
	Cout=> Carry( 	1822	),
	S=> E(	1793	));
			
  U1823	: Somador_Exato_1 PORT MAP(
	A=> C(	1887	),
	B=>E(	1732	),
	Cin=> Carry( 	1822	),
	Cout=> Carry( 	1823	),
	S=> E(	1794	));
			
  U1824	: Somador_Exato_1 PORT MAP(
	A=> C(	1888	),
	B=>E(	1733	),
	Cin=> Carry( 	1823	),
	Cout=> Carry( 	1824	),
	S=> E(	1795	));
			
  U1825	: Somador_Exato_1 PORT MAP(
	A=> C(	1889	),
	B=>E(	1734	),
	Cin=> Carry( 	1824	),
	Cout=> Carry( 	1825	),
	S=> E(	1796	));
			
  U1826	: Somador_Exato_1 PORT MAP(
	A=> C(	1890	),
	B=>E(	1735	),
	Cin=> Carry( 	1825	),
	Cout=> Carry( 	1826	),
	S=> E(	1797	));
			
  U1827	: Somador_Exato_1 PORT MAP(
	A=> C(	1891	),
	B=>E(	1736	),
	Cin=> Carry( 	1826	),
	Cout=> Carry( 	1827	),
	S=> E(	1798	));
			
  U1828	: Somador_Exato_1 PORT MAP(
	A=> C(	1892	),
	B=>E(	1737	),
	Cin=> Carry( 	1827	),
	Cout=> Carry( 	1828	),
	S=> E(	1799	));
			
  U1829	: Somador_Exato_1 PORT MAP(
	A=> C(	1893	),
	B=>E(	1738	),
	Cin=> Carry( 	1828	),
	Cout=> Carry( 	1829	),
	S=> E(	1800	));
			
  U1830	: Somador_Exato_1 PORT MAP(
	A=> C(	1894	),
	B=>E(	1739	),
	Cin=> Carry( 	1829	),
	Cout=> Carry( 	1830	),
	S=> E(	1801	));
			
  U1831	: Somador_Exato_1 PORT MAP(
	A=> C(	1895	),
	B=>E(	1740	),
	Cin=> Carry( 	1830	),
	Cout=> Carry( 	1831	),
	S=> E(	1802	));
			
  U1832	: Somador_Exato_1 PORT MAP(
	A=> C(	1896	),
	B=>E(	1741	),
	Cin=> Carry( 	1831	),
	Cout=> Carry( 	1832	),
	S=> E(	1803	));
			
  U1833	: Somador_Exato_1 PORT MAP(
	A=> C(	1897	),
	B=>E(	1742	),
	Cin=> Carry( 	1832	),
	Cout=> Carry( 	1833	),
	S=> E(	1804	));
			
  U1834	: Somador_Exato_1 PORT MAP(
	A=> C(	1898	),
	B=>E(	1743	),
	Cin=> Carry( 	1833	),
	Cout=> Carry( 	1834	),
	S=> E(	1805	));
			
  U1835	: Somador_Exato_1 PORT MAP(
	A=> C(	1899	),
	B=>E(	1744	),
	Cin=> Carry( 	1834	),
	Cout=> Carry( 	1835	),
	S=> E(	1806	));
			
  U1836	: Somador_Exato_1 PORT MAP(
	A=> C(	1900	),
	B=>E(	1745	),
	Cin=> Carry( 	1835	),
	Cout=> Carry( 	1836	),
	S=> E(	1807	));
			
  U1837	: Somador_Exato_1 PORT MAP(
	A=> C(	1901	),
	B=>E(	1746	),
	Cin=> Carry( 	1836	),
	Cout=> Carry( 	1837	),
	S=> E(	1808	));
			
  U1838	: Somador_Exato_1 PORT MAP(
	A=> C(	1902	),
	B=>E(	1747	),
	Cin=> Carry( 	1837	),
	Cout=> Carry( 	1838	),
	S=> E(	1809	));
			
  U1839	: Somador_Exato_1 PORT MAP(
	A=> C(	1903	),
	B=>E(	1748	),
	Cin=> Carry( 	1838	),
	Cout=> Carry( 	1839	),
	S=> E(	1810	));
			
  U1840	: Somador_Exato_1 PORT MAP(
	A=> C(	1904	),
	B=>E(	1749	),
	Cin=> Carry( 	1839	),
	Cout=> Carry( 	1840	),
	S=> E(	1811	));
			
  U1841	: Somador_Exato_1 PORT MAP(
	A=> C(	1905	),
	B=>E(	1750	),
	Cin=> Carry( 	1840	),
	Cout=> Carry( 	1841	),
	S=> E(	1812	));
			
  U1842	: Somador_Exato_1 PORT MAP(
	A=> C(	1906	),
	B=>E(	1751	),
	Cin=> Carry( 	1841	),
	Cout=> Carry( 	1842	),
	S=> E(	1813	));
			
  U1843	: Somador_Exato_1 PORT MAP(
	A=> C(	1907	),
	B=>E(	1752	),
	Cin=> Carry( 	1842	),
	Cout=> Carry( 	1843	),
	S=> E(	1814	));
			
  U1844	: Somador_Exato_1 PORT MAP(
	A=> C(	1908	),
	B=>E(	1753	),
	Cin=> Carry( 	1843	),
	Cout=> Carry( 	1844	),
	S=> E(	1815	));
			
  U1845	: Somador_Exato_1 PORT MAP(
	A=> C(	1909	),
	B=>E(	1754	),
	Cin=> Carry( 	1844	),
	Cout=> Carry( 	1845	),
	S=> E(	1816	));
			
  U1846	: Somador_Exato_1 PORT MAP(
	A=> C(	1910	),
	B=>E(	1755	),
	Cin=> Carry( 	1845	),
	Cout=> Carry( 	1846	),
	S=> E(	1817	));
			
  U1847	: Somador_Exato_1 PORT MAP(
	A=> C(	1911	),
	B=>E(	1756	),
	Cin=> Carry( 	1846	),
	Cout=> Carry( 	1847	),
	S=> E(	1818	));
			
  U1848	: Somador_Exato_1 PORT MAP(
	A=> C(	1912	),
	B=>E(	1757	),
	Cin=> Carry( 	1847	),
	Cout=> Carry( 	1848	),
	S=> E(	1819	));
			
  U1849	: Somador_Exato_1 PORT MAP(
	A=> C(	1913	),
	B=>E(	1758	),
	Cin=> Carry( 	1848	),
	Cout=> Carry( 	1849	),
	S=> E(	1820	));
			
  U1850	: Somador_Exato_1 PORT MAP(
	A=> C(	1914	),
	B=>E(	1759	),
	Cin=> Carry( 	1849	),
	Cout=> Carry( 	1850	),
	S=> E(	1821	));
			
  U1851	: Somador_Exato_1 PORT MAP(
	A=> C(	1915	),
	B=>E(	1760	),
	Cin=> Carry( 	1850	),
	Cout=> Carry( 	1851	),
	S=> E(	1822	));
			
  U1852	: Somador_Exato_1 PORT MAP(
	A=> C(	1916	),
	B=>E(	1761	),
	Cin=> Carry( 	1851	),
	Cout=> Carry( 	1852	),
	S=> E(	1823	));
			
  U1853	: Somador_Exato_1 PORT MAP(
	A=> C(	1917	),
	B=>E(	1762	),
	Cin=> Carry( 	1852	),
	Cout=> Carry( 	1853	),
	S=> E(	1824	));
			
  U1854	: Somador_Exato_1 PORT MAP(
	A=> C(	1918	),
	B=>E(	1763	),
	Cin=> Carry( 	1853	),
	Cout=> Carry( 	1854	),
	S=> E(	1825	));
			
  U1855	: Somador_Exato_1 PORT MAP(
	A=> C(	1919	),
	B=>Carry(	1791	),
	Cin=> Carry( 	1854	),
	Cout=> Carry( 	1855	),
	S=> E(	1826	));

			
  U1856	: Somador_Exato_1 PORT MAP(
	A=> C(	1920	),
	B=>E(	1764	),
	Cin=> '0'	,
	Cout=> Carry( 	1856	),
	S=> R(	30	));
			
  U1857	: Somador_Exato_1 PORT MAP(
	A=> C(	1921	),
	B=>E(	1765	),
	Cin=> Carry( 	1856	),
	Cout=> Carry( 	1857	),
	S=> E(	1827	));
			
  U1858	: Somador_Exato_1 PORT MAP(
	A=> C(	1922	),
	B=>E(	1766	),
	Cin=> Carry( 	1857	),
	Cout=> Carry( 	1858	),
	S=> E(	1828	));
			
  U1859	: Somador_Exato_1 PORT MAP(
	A=> C(	1923	),
	B=>E(	1767	),
	Cin=> Carry( 	1858	),
	Cout=> Carry( 	1859	),
	S=> E(	1829	));
			
  U1860	: Somador_Exato_1 PORT MAP(
	A=> C(	1924	),
	B=>E(	1768	),
	Cin=> Carry( 	1859	),
	Cout=> Carry( 	1860	),
	S=> E(	1830	));
			
  U1861	: Somador_Exato_1 PORT MAP(
	A=> C(	1925	),
	B=>E(	1769	),
	Cin=> Carry( 	1860	),
	Cout=> Carry( 	1861	),
	S=> E(	1831	));
			
  U1862	: Somador_Exato_1 PORT MAP(
	A=> C(	1926	),
	B=>E(	1770	),
	Cin=> Carry( 	1861	),
	Cout=> Carry( 	1862	),
	S=> E(	1832	));
			
  U1863	: Somador_Exato_1 PORT MAP(
	A=> C(	1927	),
	B=>E(	1771	),
	Cin=> Carry( 	1862	),
	Cout=> Carry( 	1863	),
	S=> E(	1833	));
			
  U1864	: Somador_Exato_1 PORT MAP(
	A=> C(	1928	),
	B=>E(	1772	),
	Cin=> Carry( 	1863	),
	Cout=> Carry( 	1864	),
	S=> E(	1834	));
			
  U1865	: Somador_Exato_1 PORT MAP(
	A=> C(	1929	),
	B=>E(	1773	),
	Cin=> Carry( 	1864	),
	Cout=> Carry( 	1865	),
	S=> E(	1835	));
			
  U1866	: Somador_Exato_1 PORT MAP(
	A=> C(	1930	),
	B=>E(	1774	),
	Cin=> Carry( 	1865	),
	Cout=> Carry( 	1866	),
	S=> E(	1836	));
			
  U1867	: Somador_Exato_1 PORT MAP(
	A=> C(	1931	),
	B=>E(	1775	),
	Cin=> Carry( 	1866	),
	Cout=> Carry( 	1867	),
	S=> E(	1837	));
			
  U1868	: Somador_Exato_1 PORT MAP(
	A=> C(	1932	),
	B=>E(	1776	),
	Cin=> Carry( 	1867	),
	Cout=> Carry( 	1868	),
	S=> E(	1838	));
			
  U1869	: Somador_Exato_1 PORT MAP(
	A=> C(	1933	),
	B=>E(	1777	),
	Cin=> Carry( 	1868	),
	Cout=> Carry( 	1869	),
	S=> E(	1839	));
			
  U1870	: Somador_Exato_1 PORT MAP(
	A=> C(	1934	),
	B=>E(	1778	),
	Cin=> Carry( 	1869	),
	Cout=> Carry( 	1870	),
	S=> E(	1840	));
			
  U1871	: Somador_Exato_1 PORT MAP(
	A=> C(	1935	),
	B=>E(	1779	),
	Cin=> Carry( 	1870	),
	Cout=> Carry( 	1871	),
	S=> E(	1841	));
			
  U1872	: Somador_Exato_1 PORT MAP(
	A=> C(	1936	),
	B=>E(	1780	),
	Cin=> Carry( 	1871	),
	Cout=> Carry( 	1872	),
	S=> E(	1842	));
			
  U1873	: Somador_Exato_1 PORT MAP(
	A=> C(	1937	),
	B=>E(	1781	),
	Cin=> Carry( 	1872	),
	Cout=> Carry( 	1873	),
	S=> E(	1843	));
			
  U1874	: Somador_Exato_1 PORT MAP(
	A=> C(	1938	),
	B=>E(	1782	),
	Cin=> Carry( 	1873	),
	Cout=> Carry( 	1874	),
	S=> E(	1844	));
			
  U1875	: Somador_Exato_1 PORT MAP(
	A=> C(	1939	),
	B=>E(	1783	),
	Cin=> Carry( 	1874	),
	Cout=> Carry( 	1875	),
	S=> E(	1845	));
			
  U1876	: Somador_Exato_1 PORT MAP(
	A=> C(	1940	),
	B=>E(	1784	),
	Cin=> Carry( 	1875	),
	Cout=> Carry( 	1876	),
	S=> E(	1846	));
			
  U1877	: Somador_Exato_1 PORT MAP(
	A=> C(	1941	),
	B=>E(	1785	),
	Cin=> Carry( 	1876	),
	Cout=> Carry( 	1877	),
	S=> E(	1847	));
			
  U1878	: Somador_Exato_1 PORT MAP(
	A=> C(	1942	),
	B=>E(	1786	),
	Cin=> Carry( 	1877	),
	Cout=> Carry( 	1878	),
	S=> E(	1848	));
			
  U1879	: Somador_Exato_1 PORT MAP(
	A=> C(	1943	),
	B=>E(	1787	),
	Cin=> Carry( 	1878	),
	Cout=> Carry( 	1879	),
	S=> E(	1849	));
			
  U1880	: Somador_Exato_1 PORT MAP(
	A=> C(	1944	),
	B=>E(	1788	),
	Cin=> Carry( 	1879	),
	Cout=> Carry( 	1880	),
	S=> E(	1850	));
			
  U1881	: Somador_Exato_1 PORT MAP(
	A=> C(	1945	),
	B=>E(	1789	),
	Cin=> Carry( 	1880	),
	Cout=> Carry( 	1881	),
	S=> E(	1851	));
			
  U1882	: Somador_Exato_1 PORT MAP(
	A=> C(	1946	),
	B=>E(	1790	),
	Cin=> Carry( 	1881	),
	Cout=> Carry( 	1882	),
	S=> E(	1852	));
			
  U1883	: Somador_Exato_1 PORT MAP(
	A=> C(	1947	),
	B=>E(	1791	),
	Cin=> Carry( 	1882	),
	Cout=> Carry( 	1883	),
	S=> E(	1853	));
			
  U1884	: Somador_Exato_1 PORT MAP(
	A=> C(	1948	),
	B=>E(	1792	),
	Cin=> Carry( 	1883	),
	Cout=> Carry( 	1884	),
	S=> E(	1854	));
			
  U1885	: Somador_Exato_1 PORT MAP(
	A=> C(	1949	),
	B=>E(	1793	),
	Cin=> Carry( 	1884	),
	Cout=> Carry( 	1885	),
	S=> E(	1855	));
			
  U1886	: Somador_Exato_1 PORT MAP(
	A=> C(	1950	),
	B=>E(	1794	),
	Cin=> Carry( 	1885	),
	Cout=> Carry( 	1886	),
	S=> E(	1856	));
			
  U1887	: Somador_Exato_1 PORT MAP(
	A=> C(	1951	),
	B=>E(	1795	),
	Cin=> Carry( 	1886	),
	Cout=> Carry( 	1887	),
	S=> E(	1857	));
			
  U1888	: Somador_Exato_1 PORT MAP(
	A=> C(	1952	),
	B=>E(	1796	),
	Cin=> Carry( 	1887	),
	Cout=> Carry( 	1888	),
	S=> E(	1858	));
			
  U1889	: Somador_Exato_1 PORT MAP(
	A=> C(	1953	),
	B=>E(	1797	),
	Cin=> Carry( 	1888	),
	Cout=> Carry( 	1889	),
	S=> E(	1859	));
			
  U1890	: Somador_Exato_1 PORT MAP(
	A=> C(	1954	),
	B=>E(	1798	),
	Cin=> Carry( 	1889	),
	Cout=> Carry( 	1890	),
	S=> E(	1860	));
			
  U1891	: Somador_Exato_1 PORT MAP(
	A=> C(	1955	),
	B=>E(	1799	),
	Cin=> Carry( 	1890	),
	Cout=> Carry( 	1891	),
	S=> E(	1861	));
			
  U1892	: Somador_Exato_1 PORT MAP(
	A=> C(	1956	),
	B=>E(	1800	),
	Cin=> Carry( 	1891	),
	Cout=> Carry( 	1892	),
	S=> E(	1862	));
			
  U1893	: Somador_Exato_1 PORT MAP(
	A=> C(	1957	),
	B=>E(	1801	),
	Cin=> Carry( 	1892	),
	Cout=> Carry( 	1893	),
	S=> E(	1863	));
			
  U1894	: Somador_Exato_1 PORT MAP(
	A=> C(	1958	),
	B=>E(	1802	),
	Cin=> Carry( 	1893	),
	Cout=> Carry( 	1894	),
	S=> E(	1864	));
			
  U1895	: Somador_Exato_1 PORT MAP(
	A=> C(	1959	),
	B=>E(	1803	),
	Cin=> Carry( 	1894	),
	Cout=> Carry( 	1895	),
	S=> E(	1865	));
			
  U1896	: Somador_Exato_1 PORT MAP(
	A=> C(	1960	),
	B=>E(	1804	),
	Cin=> Carry( 	1895	),
	Cout=> Carry( 	1896	),
	S=> E(	1866	));
			
  U1897	: Somador_Exato_1 PORT MAP(
	A=> C(	1961	),
	B=>E(	1805	),
	Cin=> Carry( 	1896	),
	Cout=> Carry( 	1897	),
	S=> E(	1867	));
			
  U1898	: Somador_Exato_1 PORT MAP(
	A=> C(	1962	),
	B=>E(	1806	),
	Cin=> Carry( 	1897	),
	Cout=> Carry( 	1898	),
	S=> E(	1868	));
			
  U1899	: Somador_Exato_1 PORT MAP(
	A=> C(	1963	),
	B=>E(	1807	),
	Cin=> Carry( 	1898	),
	Cout=> Carry( 	1899	),
	S=> E(	1869	));
			
  U1900	: Somador_Exato_1 PORT MAP(
	A=> C(	1964	),
	B=>E(	1808	),
	Cin=> Carry( 	1899	),
	Cout=> Carry( 	1900	),
	S=> E(	1870	));
			
  U1901	: Somador_Exato_1 PORT MAP(
	A=> C(	1965	),
	B=>E(	1809	),
	Cin=> Carry( 	1900	),
	Cout=> Carry( 	1901	),
	S=> E(	1871	));
			
  U1902	: Somador_Exato_1 PORT MAP(
	A=> C(	1966	),
	B=>E(	1810	),
	Cin=> Carry( 	1901	),
	Cout=> Carry( 	1902	),
	S=> E(	1872	));
			
  U1903	: Somador_Exato_1 PORT MAP(
	A=> C(	1967	),
	B=>E(	1811	),
	Cin=> Carry( 	1902	),
	Cout=> Carry( 	1903	),
	S=> E(	1873	));
			
  U1904	: Somador_Exato_1 PORT MAP(
	A=> C(	1968	),
	B=>E(	1812	),
	Cin=> Carry( 	1903	),
	Cout=> Carry( 	1904	),
	S=> E(	1874	));
			
  U1905	: Somador_Exato_1 PORT MAP(
	A=> C(	1969	),
	B=>E(	1813	),
	Cin=> Carry( 	1904	),
	Cout=> Carry( 	1905	),
	S=> E(	1875	));
			
  U1906	: Somador_Exato_1 PORT MAP(
	A=> C(	1970	),
	B=>E(	1814	),
	Cin=> Carry( 	1905	),
	Cout=> Carry( 	1906	),
	S=> E(	1876	));
			
  U1907	: Somador_Exato_1 PORT MAP(
	A=> C(	1971	),
	B=>E(	1815	),
	Cin=> Carry( 	1906	),
	Cout=> Carry( 	1907	),
	S=> E(	1877	));
			
  U1908	: Somador_Exato_1 PORT MAP(
	A=> C(	1972	),
	B=>E(	1816	),
	Cin=> Carry( 	1907	),
	Cout=> Carry( 	1908	),
	S=> E(	1878	));
			
  U1909	: Somador_Exato_1 PORT MAP(
	A=> C(	1973	),
	B=>E(	1817	),
	Cin=> Carry( 	1908	),
	Cout=> Carry( 	1909	),
	S=> E(	1879	));
			
  U1910	: Somador_Exato_1 PORT MAP(
	A=> C(	1974	),
	B=>E(	1818	),
	Cin=> Carry( 	1909	),
	Cout=> Carry( 	1910	),
	S=> E(	1880	));
			
  U1911	: Somador_Exato_1 PORT MAP(
	A=> C(	1975	),
	B=>E(	1819	),
	Cin=> Carry( 	1910	),
	Cout=> Carry( 	1911	),
	S=> E(	1881	));
			
  U1912	: Somador_Exato_1 PORT MAP(
	A=> C(	1976	),
	B=>E(	1820	),
	Cin=> Carry( 	1911	),
	Cout=> Carry( 	1912	),
	S=> E(	1882	));
			
  U1913	: Somador_Exato_1 PORT MAP(
	A=> C(	1977	),
	B=>E(	1821	),
	Cin=> Carry( 	1912	),
	Cout=> Carry( 	1913	),
	S=> E(	1883	));
			
  U1914	: Somador_Exato_1 PORT MAP(
	A=> C(	1978	),
	B=>E(	1822	),
	Cin=> Carry( 	1913	),
	Cout=> Carry( 	1914	),
	S=> E(	1884	));
			
  U1915	: Somador_Exato_1 PORT MAP(
	A=> C(	1979	),
	B=>E(	1823	),
	Cin=> Carry( 	1914	),
	Cout=> Carry( 	1915	),
	S=> E(	1885	));
			
  U1916	: Somador_Exato_1 PORT MAP(
	A=> C(	1980	),
	B=>E(	1824	),
	Cin=> Carry( 	1915	),
	Cout=> Carry( 	1916	),
	S=> E(	1886	));
			
  U1917	: Somador_Exato_1 PORT MAP(
	A=> C(	1981	),
	B=>E(	1825	),
	Cin=> Carry( 	1916	),
	Cout=> Carry( 	1917	),
	S=> E(	1887	));
			
  U1918	: Somador_Exato_1 PORT MAP(
	A=> C(	1982	),
	B=>E(	1826	),
	Cin=> Carry( 	1917	),
	Cout=> Carry( 	1918	),
	S=> E(	1888	));
			
  U1919	: Somador_Exato_1 PORT MAP(
	A=> C(	1983	),
	B=>Carry(	1855	),
	Cin=> Carry( 	1918	),
	Cout=> Carry( 	1919	),
	S=> E(	1889	));

			
  U1920	: Somador_Exato_1 PORT MAP(
	A=> C(	1984	),
	B=>E(	1827	),
	Cin=> '0'	,
	Cout=> Carry( 	1920	),
	S=> R(	31	));
			
  U1921	: Somador_Exato_1 PORT MAP(
	A=> C(	1985	),
	B=>E(	1828	),
	Cin=> Carry( 	1920	),
	Cout=> Carry( 	1921	),
	S=> E(	1890	));
			
  U1922	: Somador_Exato_1 PORT MAP(
	A=> C(	1986	),
	B=>E(	1829	),
	Cin=> Carry( 	1921	),
	Cout=> Carry( 	1922	),
	S=> E(	1891	));
			
  U1923	: Somador_Exato_1 PORT MAP(
	A=> C(	1987	),
	B=>E(	1830	),
	Cin=> Carry( 	1922	),
	Cout=> Carry( 	1923	),
	S=> E(	1892	));
			
  U1924	: Somador_Exato_1 PORT MAP(
	A=> C(	1988	),
	B=>E(	1831	),
	Cin=> Carry( 	1923	),
	Cout=> Carry( 	1924	),
	S=> E(	1893	));
			
  U1925	: Somador_Exato_1 PORT MAP(
	A=> C(	1989	),
	B=>E(	1832	),
	Cin=> Carry( 	1924	),
	Cout=> Carry( 	1925	),
	S=> E(	1894	));
			
  U1926	: Somador_Exato_1 PORT MAP(
	A=> C(	1990	),
	B=>E(	1833	),
	Cin=> Carry( 	1925	),
	Cout=> Carry( 	1926	),
	S=> E(	1895	));
			
  U1927	: Somador_Exato_1 PORT MAP(
	A=> C(	1991	),
	B=>E(	1834	),
	Cin=> Carry( 	1926	),
	Cout=> Carry( 	1927	),
	S=> E(	1896	));
			
  U1928	: Somador_Exato_1 PORT MAP(
	A=> C(	1992	),
	B=>E(	1835	),
	Cin=> Carry( 	1927	),
	Cout=> Carry( 	1928	),
	S=> E(	1897	));
			
  U1929	: Somador_Exato_1 PORT MAP(
	A=> C(	1993	),
	B=>E(	1836	),
	Cin=> Carry( 	1928	),
	Cout=> Carry( 	1929	),
	S=> E(	1898	));
			
  U1930	: Somador_Exato_1 PORT MAP(
	A=> C(	1994	),
	B=>E(	1837	),
	Cin=> Carry( 	1929	),
	Cout=> Carry( 	1930	),
	S=> E(	1899	));
			
  U1931	: Somador_Exato_1 PORT MAP(
	A=> C(	1995	),
	B=>E(	1838	),
	Cin=> Carry( 	1930	),
	Cout=> Carry( 	1931	),
	S=> E(	1900	));
			
  U1932	: Somador_Exato_1 PORT MAP(
	A=> C(	1996	),
	B=>E(	1839	),
	Cin=> Carry( 	1931	),
	Cout=> Carry( 	1932	),
	S=> E(	1901	));
			
  U1933	: Somador_Exato_1 PORT MAP(
	A=> C(	1997	),
	B=>E(	1840	),
	Cin=> Carry( 	1932	),
	Cout=> Carry( 	1933	),
	S=> E(	1902	));
			
  U1934	: Somador_Exato_1 PORT MAP(
	A=> C(	1998	),
	B=>E(	1841	),
	Cin=> Carry( 	1933	),
	Cout=> Carry( 	1934	),
	S=> E(	1903	));
			
  U1935	: Somador_Exato_1 PORT MAP(
	A=> C(	1999	),
	B=>E(	1842	),
	Cin=> Carry( 	1934	),
	Cout=> Carry( 	1935	),
	S=> E(	1904	));
			
  U1936	: Somador_Exato_1 PORT MAP(
	A=> C(	2000	),
	B=>E(	1843	),
	Cin=> Carry( 	1935	),
	Cout=> Carry( 	1936	),
	S=> E(	1905	));
			
  U1937	: Somador_Exato_1 PORT MAP(
	A=> C(	2001	),
	B=>E(	1844	),
	Cin=> Carry( 	1936	),
	Cout=> Carry( 	1937	),
	S=> E(	1906	));
			
  U1938	: Somador_Exato_1 PORT MAP(
	A=> C(	2002	),
	B=>E(	1845	),
	Cin=> Carry( 	1937	),
	Cout=> Carry( 	1938	),
	S=> E(	1907	));
			
  U1939	: Somador_Exato_1 PORT MAP(
	A=> C(	2003	),
	B=>E(	1846	),
	Cin=> Carry( 	1938	),
	Cout=> Carry( 	1939	),
	S=> E(	1908	));
			
  U1940	: Somador_Exato_1 PORT MAP(
	A=> C(	2004	),
	B=>E(	1847	),
	Cin=> Carry( 	1939	),
	Cout=> Carry( 	1940	),
	S=> E(	1909	));
			
  U1941	: Somador_Exato_1 PORT MAP(
	A=> C(	2005	),
	B=>E(	1848	),
	Cin=> Carry( 	1940	),
	Cout=> Carry( 	1941	),
	S=> E(	1910	));
			
  U1942	: Somador_Exato_1 PORT MAP(
	A=> C(	2006	),
	B=>E(	1849	),
	Cin=> Carry( 	1941	),
	Cout=> Carry( 	1942	),
	S=> E(	1911	));
			
  U1943	: Somador_Exato_1 PORT MAP(
	A=> C(	2007	),
	B=>E(	1850	),
	Cin=> Carry( 	1942	),
	Cout=> Carry( 	1943	),
	S=> E(	1912	));
			
  U1944	: Somador_Exato_1 PORT MAP(
	A=> C(	2008	),
	B=>E(	1851	),
	Cin=> Carry( 	1943	),
	Cout=> Carry( 	1944	),
	S=> E(	1913	));
			
  U1945	: Somador_Exato_1 PORT MAP(
	A=> C(	2009	),
	B=>E(	1852	),
	Cin=> Carry( 	1944	),
	Cout=> Carry( 	1945	),
	S=> E(	1914	));
			
  U1946	: Somador_Exato_1 PORT MAP(
	A=> C(	2010	),
	B=>E(	1853	),
	Cin=> Carry( 	1945	),
	Cout=> Carry( 	1946	),
	S=> E(	1915	));
			
  U1947	: Somador_Exato_1 PORT MAP(
	A=> C(	2011	),
	B=>E(	1854	),
	Cin=> Carry( 	1946	),
	Cout=> Carry( 	1947	),
	S=> E(	1916	));
			
  U1948	: Somador_Exato_1 PORT MAP(
	A=> C(	2012	),
	B=>E(	1855	),
	Cin=> Carry( 	1947	),
	Cout=> Carry( 	1948	),
	S=> E(	1917	));
			
  U1949	: Somador_Exato_1 PORT MAP(
	A=> C(	2013	),
	B=>E(	1856	),
	Cin=> Carry( 	1948	),
	Cout=> Carry( 	1949	),
	S=> E(	1918	));
			
  U1950	: Somador_Exato_1 PORT MAP(
	A=> C(	2014	),
	B=>E(	1857	),
	Cin=> Carry( 	1949	),
	Cout=> Carry( 	1950	),
	S=> E(	1919	));
			
  U1951	: Somador_Exato_1 PORT MAP(
	A=> C(	2015	),
	B=>E(	1858	),
	Cin=> Carry( 	1950	),
	Cout=> Carry( 	1951	),
	S=> E(	1920	));
			
  U1952	: Somador_Exato_1 PORT MAP(
	A=> C(	2016	),
	B=>E(	1859	),
	Cin=> Carry( 	1951	),
	Cout=> Carry( 	1952	),
	S=> E(	1921	));
			
  U1953	: Somador_Exato_1 PORT MAP(
	A=> C(	2017	),
	B=>E(	1860	),
	Cin=> Carry( 	1952	),
	Cout=> Carry( 	1953	),
	S=> E(	1922	));
			
  U1954	: Somador_Exato_1 PORT MAP(
	A=> C(	2018	),
	B=>E(	1861	),
	Cin=> Carry( 	1953	),
	Cout=> Carry( 	1954	),
	S=> E(	1923	));
			
  U1955	: Somador_Exato_1 PORT MAP(
	A=> C(	2019	),
	B=>E(	1862	),
	Cin=> Carry( 	1954	),
	Cout=> Carry( 	1955	),
	S=> E(	1924	));
			
  U1956	: Somador_Exato_1 PORT MAP(
	A=> C(	2020	),
	B=>E(	1863	),
	Cin=> Carry( 	1955	),
	Cout=> Carry( 	1956	),
	S=> E(	1925	));
			
  U1957	: Somador_Exato_1 PORT MAP(
	A=> C(	2021	),
	B=>E(	1864	),
	Cin=> Carry( 	1956	),
	Cout=> Carry( 	1957	),
	S=> E(	1926	));
			
  U1958	: Somador_Exato_1 PORT MAP(
	A=> C(	2022	),
	B=>E(	1865	),
	Cin=> Carry( 	1957	),
	Cout=> Carry( 	1958	),
	S=> E(	1927	));
			
  U1959	: Somador_Exato_1 PORT MAP(
	A=> C(	2023	),
	B=>E(	1866	),
	Cin=> Carry( 	1958	),
	Cout=> Carry( 	1959	),
	S=> E(	1928	));
			
  U1960	: Somador_Exato_1 PORT MAP(
	A=> C(	2024	),
	B=>E(	1867	),
	Cin=> Carry( 	1959	),
	Cout=> Carry( 	1960	),
	S=> E(	1929	));
			
  U1961	: Somador_Exato_1 PORT MAP(
	A=> C(	2025	),
	B=>E(	1868	),
	Cin=> Carry( 	1960	),
	Cout=> Carry( 	1961	),
	S=> E(	1930	));
			
  U1962	: Somador_Exato_1 PORT MAP(
	A=> C(	2026	),
	B=>E(	1869	),
	Cin=> Carry( 	1961	),
	Cout=> Carry( 	1962	),
	S=> E(	1931	));
			
  U1963	: Somador_Exato_1 PORT MAP(
	A=> C(	2027	),
	B=>E(	1870	),
	Cin=> Carry( 	1962	),
	Cout=> Carry( 	1963	),
	S=> E(	1932	));
			
  U1964	: Somador_Exato_1 PORT MAP(
	A=> C(	2028	),
	B=>E(	1871	),
	Cin=> Carry( 	1963	),
	Cout=> Carry( 	1964	),
	S=> E(	1933	));
			
  U1965	: Somador_Exato_1 PORT MAP(
	A=> C(	2029	),
	B=>E(	1872	),
	Cin=> Carry( 	1964	),
	Cout=> Carry( 	1965	),
	S=> E(	1934	));
			
  U1966	: Somador_Exato_1 PORT MAP(
	A=> C(	2030	),
	B=>E(	1873	),
	Cin=> Carry( 	1965	),
	Cout=> Carry( 	1966	),
	S=> E(	1935	));
			
  U1967	: Somador_Exato_1 PORT MAP(
	A=> C(	2031	),
	B=>E(	1874	),
	Cin=> Carry( 	1966	),
	Cout=> Carry( 	1967	),
	S=> E(	1936	));
			
  U1968	: Somador_Exato_1 PORT MAP(
	A=> C(	2032	),
	B=>E(	1875	),
	Cin=> Carry( 	1967	),
	Cout=> Carry( 	1968	),
	S=> E(	1937	));
			
  U1969	: Somador_Exato_1 PORT MAP(
	A=> C(	2033	),
	B=>E(	1876	),
	Cin=> Carry( 	1968	),
	Cout=> Carry( 	1969	),
	S=> E(	1938	));
			
  U1970	: Somador_Exato_1 PORT MAP(
	A=> C(	2034	),
	B=>E(	1877	),
	Cin=> Carry( 	1969	),
	Cout=> Carry( 	1970	),
	S=> E(	1939	));
			
  U1971	: Somador_Exato_1 PORT MAP(
	A=> C(	2035	),
	B=>E(	1878	),
	Cin=> Carry( 	1970	),
	Cout=> Carry( 	1971	),
	S=> E(	1940	));
			
  U1972	: Somador_Exato_1 PORT MAP(
	A=> C(	2036	),
	B=>E(	1879	),
	Cin=> Carry( 	1971	),
	Cout=> Carry( 	1972	),
	S=> E(	1941	));
			
  U1973	: Somador_Exato_1 PORT MAP(
	A=> C(	2037	),
	B=>E(	1880	),
	Cin=> Carry( 	1972	),
	Cout=> Carry( 	1973	),
	S=> E(	1942	));
			
  U1974	: Somador_Exato_1 PORT MAP(
	A=> C(	2038	),
	B=>E(	1881	),
	Cin=> Carry( 	1973	),
	Cout=> Carry( 	1974	),
	S=> E(	1943	));
			
  U1975	: Somador_Exato_1 PORT MAP(
	A=> C(	2039	),
	B=>E(	1882	),
	Cin=> Carry( 	1974	),
	Cout=> Carry( 	1975	),
	S=> E(	1944	));
			
  U1976	: Somador_Exato_1 PORT MAP(
	A=> C(	2040	),
	B=>E(	1883	),
	Cin=> Carry( 	1975	),
	Cout=> Carry( 	1976	),
	S=> E(	1945	));
			
  U1977	: Somador_Exato_1 PORT MAP(
	A=> C(	2041	),
	B=>E(	1884	),
	Cin=> Carry( 	1976	),
	Cout=> Carry( 	1977	),
	S=> E(	1946	));
			
  U1978	: Somador_Exato_1 PORT MAP(
	A=> C(	2042	),
	B=>E(	1885	),
	Cin=> Carry( 	1977	),
	Cout=> Carry( 	1978	),
	S=> E(	1947	));
			
  U1979	: Somador_Exato_1 PORT MAP(
	A=> C(	2043	),
	B=>E(	1886	),
	Cin=> Carry( 	1978	),
	Cout=> Carry( 	1979	),
	S=> E(	1948	));
			
  U1980	: Somador_Exato_1 PORT MAP(
	A=> C(	2044	),
	B=>E(	1887	),
	Cin=> Carry( 	1979	),
	Cout=> Carry( 	1980	),
	S=> E(	1949	));
			
  U1981	: Somador_Exato_1 PORT MAP(
	A=> C(	2045	),
	B=>E(	1888	),
	Cin=> Carry( 	1980	),
	Cout=> Carry( 	1981	),
	S=> E(	1950	));
			
  U1982	: Somador_Exato_1 PORT MAP(
	A=> C(	2046	),
	B=>E(	1889	),
	Cin=> Carry( 	1981	),
	Cout=> Carry( 	1982	),
	S=> E(	1951	));
			
  U1983	: Somador_Exato_1 PORT MAP(
	A=> C(	2047	),
	B=>Carry(	1919	),
	Cin=> Carry( 	1982	),
	Cout=> Carry( 	1983	),
	S=> E(	1952	));

			
  U1984	: Somador_Exato_1 PORT MAP(
	A=> C(	2048	),
	B=>E(	1890	),
	Cin=> '0'	,
	Cout=> Carry( 	1984	),
	S=> R(	32	));
			
  U1985	: Somador_Exato_1 PORT MAP(
	A=> C(	2049	),
	B=>E(	1891	),
	Cin=> Carry( 	1984	),
	Cout=> Carry( 	1985	),
	S=> E(	1953	));
			
  U1986	: Somador_Exato_1 PORT MAP(
	A=> C(	2050	),
	B=>E(	1892	),
	Cin=> Carry( 	1985	),
	Cout=> Carry( 	1986	),
	S=> E(	1954	));
			
  U1987	: Somador_Exato_1 PORT MAP(
	A=> C(	2051	),
	B=>E(	1893	),
	Cin=> Carry( 	1986	),
	Cout=> Carry( 	1987	),
	S=> E(	1955	));
			
  U1988	: Somador_Exato_1 PORT MAP(
	A=> C(	2052	),
	B=>E(	1894	),
	Cin=> Carry( 	1987	),
	Cout=> Carry( 	1988	),
	S=> E(	1956	));
			
  U1989	: Somador_Exato_1 PORT MAP(
	A=> C(	2053	),
	B=>E(	1895	),
	Cin=> Carry( 	1988	),
	Cout=> Carry( 	1989	),
	S=> E(	1957	));
			
  U1990	: Somador_Exato_1 PORT MAP(
	A=> C(	2054	),
	B=>E(	1896	),
	Cin=> Carry( 	1989	),
	Cout=> Carry( 	1990	),
	S=> E(	1958	));
			
  U1991	: Somador_Exato_1 PORT MAP(
	A=> C(	2055	),
	B=>E(	1897	),
	Cin=> Carry( 	1990	),
	Cout=> Carry( 	1991	),
	S=> E(	1959	));
			
  U1992	: Somador_Exato_1 PORT MAP(
	A=> C(	2056	),
	B=>E(	1898	),
	Cin=> Carry( 	1991	),
	Cout=> Carry( 	1992	),
	S=> E(	1960	));
			
  U1993	: Somador_Exato_1 PORT MAP(
	A=> C(	2057	),
	B=>E(	1899	),
	Cin=> Carry( 	1992	),
	Cout=> Carry( 	1993	),
	S=> E(	1961	));
			
  U1994	: Somador_Exato_1 PORT MAP(
	A=> C(	2058	),
	B=>E(	1900	),
	Cin=> Carry( 	1993	),
	Cout=> Carry( 	1994	),
	S=> E(	1962	));
			
  U1995	: Somador_Exato_1 PORT MAP(
	A=> C(	2059	),
	B=>E(	1901	),
	Cin=> Carry( 	1994	),
	Cout=> Carry( 	1995	),
	S=> E(	1963	));
			
  U1996	: Somador_Exato_1 PORT MAP(
	A=> C(	2060	),
	B=>E(	1902	),
	Cin=> Carry( 	1995	),
	Cout=> Carry( 	1996	),
	S=> E(	1964	));
			
  U1997	: Somador_Exato_1 PORT MAP(
	A=> C(	2061	),
	B=>E(	1903	),
	Cin=> Carry( 	1996	),
	Cout=> Carry( 	1997	),
	S=> E(	1965	));
			
  U1998	: Somador_Exato_1 PORT MAP(
	A=> C(	2062	),
	B=>E(	1904	),
	Cin=> Carry( 	1997	),
	Cout=> Carry( 	1998	),
	S=> E(	1966	));
			
  U1999	: Somador_Exato_1 PORT MAP(
	A=> C(	2063	),
	B=>E(	1905	),
	Cin=> Carry( 	1998	),
	Cout=> Carry( 	1999	),
	S=> E(	1967	));
			
  U2000	: Somador_Exato_1 PORT MAP(
	A=> C(	2064	),
	B=>E(	1906	),
	Cin=> Carry( 	1999	),
	Cout=> Carry( 	2000	),
	S=> E(	1968	));
			
  U2001	: Somador_Exato_1 PORT MAP(
	A=> C(	2065	),
	B=>E(	1907	),
	Cin=> Carry( 	2000	),
	Cout=> Carry( 	2001	),
	S=> E(	1969	));
			
  U2002	: Somador_Exato_1 PORT MAP(
	A=> C(	2066	),
	B=>E(	1908	),
	Cin=> Carry( 	2001	),
	Cout=> Carry( 	2002	),
	S=> E(	1970	));
			
  U2003	: Somador_Exato_1 PORT MAP(
	A=> C(	2067	),
	B=>E(	1909	),
	Cin=> Carry( 	2002	),
	Cout=> Carry( 	2003	),
	S=> E(	1971	));
			
  U2004	: Somador_Exato_1 PORT MAP(
	A=> C(	2068	),
	B=>E(	1910	),
	Cin=> Carry( 	2003	),
	Cout=> Carry( 	2004	),
	S=> E(	1972	));
			
  U2005	: Somador_Exato_1 PORT MAP(
	A=> C(	2069	),
	B=>E(	1911	),
	Cin=> Carry( 	2004	),
	Cout=> Carry( 	2005	),
	S=> E(	1973	));
			
  U2006	: Somador_Exato_1 PORT MAP(
	A=> C(	2070	),
	B=>E(	1912	),
	Cin=> Carry( 	2005	),
	Cout=> Carry( 	2006	),
	S=> E(	1974	));
			
  U2007	: Somador_Exato_1 PORT MAP(
	A=> C(	2071	),
	B=>E(	1913	),
	Cin=> Carry( 	2006	),
	Cout=> Carry( 	2007	),
	S=> E(	1975	));
			
  U2008	: Somador_Exato_1 PORT MAP(
	A=> C(	2072	),
	B=>E(	1914	),
	Cin=> Carry( 	2007	),
	Cout=> Carry( 	2008	),
	S=> E(	1976	));
			
  U2009	: Somador_Exato_1 PORT MAP(
	A=> C(	2073	),
	B=>E(	1915	),
	Cin=> Carry( 	2008	),
	Cout=> Carry( 	2009	),
	S=> E(	1977	));
			
  U2010	: Somador_Exato_1 PORT MAP(
	A=> C(	2074	),
	B=>E(	1916	),
	Cin=> Carry( 	2009	),
	Cout=> Carry( 	2010	),
	S=> E(	1978	));
			
  U2011	: Somador_Exato_1 PORT MAP(
	A=> C(	2075	),
	B=>E(	1917	),
	Cin=> Carry( 	2010	),
	Cout=> Carry( 	2011	),
	S=> E(	1979	));
			
  U2012	: Somador_Exato_1 PORT MAP(
	A=> C(	2076	),
	B=>E(	1918	),
	Cin=> Carry( 	2011	),
	Cout=> Carry( 	2012	),
	S=> E(	1980	));
			
  U2013	: Somador_Exato_1 PORT MAP(
	A=> C(	2077	),
	B=>E(	1919	),
	Cin=> Carry( 	2012	),
	Cout=> Carry( 	2013	),
	S=> E(	1981	));
			
  U2014	: Somador_Exato_1 PORT MAP(
	A=> C(	2078	),
	B=>E(	1920	),
	Cin=> Carry( 	2013	),
	Cout=> Carry( 	2014	),
	S=> E(	1982	));
			
  U2015	: Somador_Exato_1 PORT MAP(
	A=> C(	2079	),
	B=>E(	1921	),
	Cin=> Carry( 	2014	),
	Cout=> Carry( 	2015	),
	S=> E(	1983	));
			
  U2016	: Soma_AMA3_1 PORT MAP(
	A=> C(	2080	),
	B=>E(	1922	),
	Cin=> Carry( 	2015	),
	Cout=> Carry( 	2016	),
	S=> E(	1984	));
			
  U2017	: Soma_AMA3_1 PORT MAP(
	A=> C(	2081	),
	B=>E(	1923	),
	Cin=> Carry( 	2016	),
	Cout=> Carry( 	2017	),
	S=> E(	1985	));
			
  U2018	: Soma_AMA3_1 PORT MAP(
	A=> C(	2082	),
	B=>E(	1924	),
	Cin=> Carry( 	2017	),
	Cout=> Carry( 	2018	),
	S=> E(	1986	));
			
  U2019	: Soma_AMA3_1 PORT MAP(
	A=> C(	2083	),
	B=>E(	1925	),
	Cin=> Carry( 	2018	),
	Cout=> Carry( 	2019	),
	S=> E(	1987	));
			
  U2020	: Soma_AMA3_1 PORT MAP(
	A=> C(	2084	),
	B=>E(	1926	),
	Cin=> Carry( 	2019	),
	Cout=> Carry( 	2020	),
	S=> E(	1988	));
			
  U2021	: Soma_AMA3_1 PORT MAP(
	A=> C(	2085	),
	B=>E(	1927	),
	Cin=> Carry( 	2020	),
	Cout=> Carry( 	2021	),
	S=> E(	1989	));
			
  U2022	: Soma_AMA3_1 PORT MAP(
	A=> C(	2086	),
	B=>E(	1928	),
	Cin=> Carry( 	2021	),
	Cout=> Carry( 	2022	),
	S=> E(	1990	));
			
  U2023	: Soma_AMA3_1 PORT MAP(
	A=> C(	2087	),
	B=>E(	1929	),
	Cin=> Carry( 	2022	),
	Cout=> Carry( 	2023	),
	S=> E(	1991	));
			
  U2024	: Soma_AMA3_1 PORT MAP(
	A=> C(	2088	),
	B=>E(	1930	),
	Cin=> Carry( 	2023	),
	Cout=> Carry( 	2024	),
	S=> E(	1992	));
			
  U2025	: Soma_AMA3_1 PORT MAP(
	A=> C(	2089	),
	B=>E(	1931	),
	Cin=> Carry( 	2024	),
	Cout=> Carry( 	2025	),
	S=> E(	1993	));
			
  U2026	: Soma_AMA3_1 PORT MAP(
	A=> C(	2090	),
	B=>E(	1932	),
	Cin=> Carry( 	2025	),
	Cout=> Carry( 	2026	),
	S=> E(	1994	));
			
  U2027	: Soma_AMA3_1 PORT MAP(
	A=> C(	2091	),
	B=>E(	1933	),
	Cin=> Carry( 	2026	),
	Cout=> Carry( 	2027	),
	S=> E(	1995	));
			
  U2028	: Soma_AMA3_1 PORT MAP(
	A=> C(	2092	),
	B=>E(	1934	),
	Cin=> Carry( 	2027	),
	Cout=> Carry( 	2028	),
	S=> E(	1996	));
			
  U2029	: Soma_AMA3_1 PORT MAP(
	A=> C(	2093	),
	B=>E(	1935	),
	Cin=> Carry( 	2028	),
	Cout=> Carry( 	2029	),
	S=> E(	1997	));
			
  U2030	: Soma_AMA3_1 PORT MAP(
	A=> C(	2094	),
	B=>E(	1936	),
	Cin=> Carry( 	2029	),
	Cout=> Carry( 	2030	),
	S=> E(	1998	));
			
  U2031	: Soma_AMA3_1 PORT MAP(
	A=> C(	2095	),
	B=>E(	1937	),
	Cin=> Carry( 	2030	),
	Cout=> Carry( 	2031	),
	S=> E(	1999	));
			
  U2032	: Soma_AMA3_1 PORT MAP(
	A=> C(	2096	),
	B=>E(	1938	),
	Cin=> Carry( 	2031	),
	Cout=> Carry( 	2032	),
	S=> E(	2000	));
			
  U2033	: Soma_AMA3_1 PORT MAP(
	A=> C(	2097	),
	B=>E(	1939	),
	Cin=> Carry( 	2032	),
	Cout=> Carry( 	2033	),
	S=> E(	2001	));
			
  U2034	: Soma_AMA3_1 PORT MAP(
	A=> C(	2098	),
	B=>E(	1940	),
	Cin=> Carry( 	2033	),
	Cout=> Carry( 	2034	),
	S=> E(	2002	));
			
  U2035	: Soma_AMA3_1 PORT MAP(
	A=> C(	2099	),
	B=>E(	1941	),
	Cin=> Carry( 	2034	),
	Cout=> Carry( 	2035	),
	S=> E(	2003	));
			
  U2036	: Soma_AMA3_1 PORT MAP(
	A=> C(	2100	),
	B=>E(	1942	),
	Cin=> Carry( 	2035	),
	Cout=> Carry( 	2036	),
	S=> E(	2004	));
			
  U2037	: Soma_AMA3_1 PORT MAP(
	A=> C(	2101	),
	B=>E(	1943	),
	Cin=> Carry( 	2036	),
	Cout=> Carry( 	2037	),
	S=> E(	2005	));
			
  U2038	: Soma_AMA3_1 PORT MAP(
	A=> C(	2102	),
	B=>E(	1944	),
	Cin=> Carry( 	2037	),
	Cout=> Carry( 	2038	),
	S=> E(	2006	));
			
  U2039	: Soma_AMA3_1 PORT MAP(
	A=> C(	2103	),
	B=>E(	1945	),
	Cin=> Carry( 	2038	),
	Cout=> Carry( 	2039	),
	S=> E(	2007	));
			
  U2040	: Soma_AMA3_1 PORT MAP(
	A=> C(	2104	),
	B=>E(	1946	),
	Cin=> Carry( 	2039	),
	Cout=> Carry( 	2040	),
	S=> E(	2008	));
			
  U2041	: Soma_AMA3_1 PORT MAP(
	A=> C(	2105	),
	B=>E(	1947	),
	Cin=> Carry( 	2040	),
	Cout=> Carry( 	2041	),
	S=> E(	2009	));
			
  U2042	: Soma_AMA3_1 PORT MAP(
	A=> C(	2106	),
	B=>E(	1948	),
	Cin=> Carry( 	2041	),
	Cout=> Carry( 	2042	),
	S=> E(	2010	));
			
  U2043	: Soma_AMA3_1 PORT MAP(
	A=> C(	2107	),
	B=>E(	1949	),
	Cin=> Carry( 	2042	),
	Cout=> Carry( 	2043	),
	S=> E(	2011	));
			
  U2044	: Soma_AMA3_1 PORT MAP(
	A=> C(	2108	),
	B=>E(	1950	),
	Cin=> Carry( 	2043	),
	Cout=> Carry( 	2044	),
	S=> E(	2012	));
			
  U2045	: Soma_AMA3_1 PORT MAP(
	A=> C(	2109	),
	B=>E(	1951	),
	Cin=> Carry( 	2044	),
	Cout=> Carry( 	2045	),
	S=> E(	2013	));
			
  U2046	: Soma_AMA3_1 PORT MAP(
	A=> C(	2110	),
	B=>E(	1952	),
	Cin=> Carry( 	2045	),
	Cout=> Carry( 	2046	),
	S=> E(	2014	));
			
  U2047	: Soma_AMA3_1 PORT MAP(
	A=> C(	2111	),
	B=>Carry(	1983	),
	Cin=> Carry( 	2046	),
	Cout=> Carry( 	2047	),
	S=> E(	2015	));

			
  U2048	: Soma_AMA3_1 PORT MAP(
	A=> C(	2112	),
	B=>E(	1953	),
	Cin=> '0'	,
	Cout=> Carry( 	2048	),
	S=> R(	33	));
			
  U2049	: Soma_AMA3_1 PORT MAP(
	A=> C(	2113	),
	B=>E(	1954	),
	Cin=> Carry( 	2048	),
	Cout=> Carry( 	2049	),
	S=> E(	2016	));
			
  U2050	: Soma_AMA3_1 PORT MAP(
	A=> C(	2114	),
	B=>E(	1955	),
	Cin=> Carry( 	2049	),
	Cout=> Carry( 	2050	),
	S=> E(	2017	));
			
  U2051	: Soma_AMA3_1 PORT MAP(
	A=> C(	2115	),
	B=>E(	1956	),
	Cin=> Carry( 	2050	),
	Cout=> Carry( 	2051	),
	S=> E(	2018	));
			
  U2052	: Soma_AMA3_1 PORT MAP(
	A=> C(	2116	),
	B=>E(	1957	),
	Cin=> Carry( 	2051	),
	Cout=> Carry( 	2052	),
	S=> E(	2019	));
			
  U2053	: Soma_AMA3_1 PORT MAP(
	A=> C(	2117	),
	B=>E(	1958	),
	Cin=> Carry( 	2052	),
	Cout=> Carry( 	2053	),
	S=> E(	2020	));
			
  U2054	: Soma_AMA3_1 PORT MAP(
	A=> C(	2118	),
	B=>E(	1959	),
	Cin=> Carry( 	2053	),
	Cout=> Carry( 	2054	),
	S=> E(	2021	));
			
  U2055	: Soma_AMA3_1 PORT MAP(
	A=> C(	2119	),
	B=>E(	1960	),
	Cin=> Carry( 	2054	),
	Cout=> Carry( 	2055	),
	S=> E(	2022	));
			
  U2056	: Soma_AMA3_1 PORT MAP(
	A=> C(	2120	),
	B=>E(	1961	),
	Cin=> Carry( 	2055	),
	Cout=> Carry( 	2056	),
	S=> E(	2023	));
			
  U2057	: Soma_AMA3_1 PORT MAP(
	A=> C(	2121	),
	B=>E(	1962	),
	Cin=> Carry( 	2056	),
	Cout=> Carry( 	2057	),
	S=> E(	2024	));
			
  U2058	: Soma_AMA3_1 PORT MAP(
	A=> C(	2122	),
	B=>E(	1963	),
	Cin=> Carry( 	2057	),
	Cout=> Carry( 	2058	),
	S=> E(	2025	));
			
  U2059	: Soma_AMA3_1 PORT MAP(
	A=> C(	2123	),
	B=>E(	1964	),
	Cin=> Carry( 	2058	),
	Cout=> Carry( 	2059	),
	S=> E(	2026	));
			
  U2060	: Soma_AMA3_1 PORT MAP(
	A=> C(	2124	),
	B=>E(	1965	),
	Cin=> Carry( 	2059	),
	Cout=> Carry( 	2060	),
	S=> E(	2027	));
			
  U2061	: Soma_AMA3_1 PORT MAP(
	A=> C(	2125	),
	B=>E(	1966	),
	Cin=> Carry( 	2060	),
	Cout=> Carry( 	2061	),
	S=> E(	2028	));
			
  U2062	: Soma_AMA3_1 PORT MAP(
	A=> C(	2126	),
	B=>E(	1967	),
	Cin=> Carry( 	2061	),
	Cout=> Carry( 	2062	),
	S=> E(	2029	));
			
  U2063	: Soma_AMA3_1 PORT MAP(
	A=> C(	2127	),
	B=>E(	1968	),
	Cin=> Carry( 	2062	),
	Cout=> Carry( 	2063	),
	S=> E(	2030	));
			
  U2064	: Soma_AMA3_1 PORT MAP(
	A=> C(	2128	),
	B=>E(	1969	),
	Cin=> Carry( 	2063	),
	Cout=> Carry( 	2064	),
	S=> E(	2031	));
			
  U2065	: Soma_AMA3_1 PORT MAP(
	A=> C(	2129	),
	B=>E(	1970	),
	Cin=> Carry( 	2064	),
	Cout=> Carry( 	2065	),
	S=> E(	2032	));
			
  U2066	: Soma_AMA3_1 PORT MAP(
	A=> C(	2130	),
	B=>E(	1971	),
	Cin=> Carry( 	2065	),
	Cout=> Carry( 	2066	),
	S=> E(	2033	));
			
  U2067	: Soma_AMA3_1 PORT MAP(
	A=> C(	2131	),
	B=>E(	1972	),
	Cin=> Carry( 	2066	),
	Cout=> Carry( 	2067	),
	S=> E(	2034	));
			
  U2068	: Soma_AMA3_1 PORT MAP(
	A=> C(	2132	),
	B=>E(	1973	),
	Cin=> Carry( 	2067	),
	Cout=> Carry( 	2068	),
	S=> E(	2035	));
			
  U2069	: Soma_AMA3_1 PORT MAP(
	A=> C(	2133	),
	B=>E(	1974	),
	Cin=> Carry( 	2068	),
	Cout=> Carry( 	2069	),
	S=> E(	2036	));
			
  U2070	: Soma_AMA3_1 PORT MAP(
	A=> C(	2134	),
	B=>E(	1975	),
	Cin=> Carry( 	2069	),
	Cout=> Carry( 	2070	),
	S=> E(	2037	));
			
  U2071	: Soma_AMA3_1 PORT MAP(
	A=> C(	2135	),
	B=>E(	1976	),
	Cin=> Carry( 	2070	),
	Cout=> Carry( 	2071	),
	S=> E(	2038	));
			
  U2072	: Soma_AMA3_1 PORT MAP(
	A=> C(	2136	),
	B=>E(	1977	),
	Cin=> Carry( 	2071	),
	Cout=> Carry( 	2072	),
	S=> E(	2039	));
			
  U2073	: Soma_AMA3_1 PORT MAP(
	A=> C(	2137	),
	B=>E(	1978	),
	Cin=> Carry( 	2072	),
	Cout=> Carry( 	2073	),
	S=> E(	2040	));
			
  U2074	: Soma_AMA3_1 PORT MAP(
	A=> C(	2138	),
	B=>E(	1979	),
	Cin=> Carry( 	2073	),
	Cout=> Carry( 	2074	),
	S=> E(	2041	));
			
  U2075	: Soma_AMA3_1 PORT MAP(
	A=> C(	2139	),
	B=>E(	1980	),
	Cin=> Carry( 	2074	),
	Cout=> Carry( 	2075	),
	S=> E(	2042	));
			
  U2076	: Soma_AMA3_1 PORT MAP(
	A=> C(	2140	),
	B=>E(	1981	),
	Cin=> Carry( 	2075	),
	Cout=> Carry( 	2076	),
	S=> E(	2043	));
			
  U2077	: Soma_AMA3_1 PORT MAP(
	A=> C(	2141	),
	B=>E(	1982	),
	Cin=> Carry( 	2076	),
	Cout=> Carry( 	2077	),
	S=> E(	2044	));
			
  U2078	: Soma_AMA3_1 PORT MAP(
	A=> C(	2142	),
	B=>E(	1983	),
	Cin=> Carry( 	2077	),
	Cout=> Carry( 	2078	),
	S=> E(	2045	));
			
  U2079	: Soma_AMA3_1 PORT MAP(
	A=> C(	2143	),
	B=>E(	1984	),
	Cin=> Carry( 	2078	),
	Cout=> Carry( 	2079	),
	S=> E(	2046	));
			
  U2080	: Soma_AMA3_1 PORT MAP(
	A=> C(	2144	),
	B=>E(	1985	),
	Cin=> Carry( 	2079	),
	Cout=> Carry( 	2080	),
	S=> E(	2047	));
			
  U2081	: Soma_AMA3_1 PORT MAP(
	A=> C(	2145	),
	B=>E(	1986	),
	Cin=> Carry( 	2080	),
	Cout=> Carry( 	2081	),
	S=> E(	2048	));
			
  U2082	: Soma_AMA3_1 PORT MAP(
	A=> C(	2146	),
	B=>E(	1987	),
	Cin=> Carry( 	2081	),
	Cout=> Carry( 	2082	),
	S=> E(	2049	));
			
  U2083	: Soma_AMA3_1 PORT MAP(
	A=> C(	2147	),
	B=>E(	1988	),
	Cin=> Carry( 	2082	),
	Cout=> Carry( 	2083	),
	S=> E(	2050	));
			
  U2084	: Soma_AMA3_1 PORT MAP(
	A=> C(	2148	),
	B=>E(	1989	),
	Cin=> Carry( 	2083	),
	Cout=> Carry( 	2084	),
	S=> E(	2051	));
			
  U2085	: Soma_AMA3_1 PORT MAP(
	A=> C(	2149	),
	B=>E(	1990	),
	Cin=> Carry( 	2084	),
	Cout=> Carry( 	2085	),
	S=> E(	2052	));
			
  U2086	: Soma_AMA3_1 PORT MAP(
	A=> C(	2150	),
	B=>E(	1991	),
	Cin=> Carry( 	2085	),
	Cout=> Carry( 	2086	),
	S=> E(	2053	));
			
  U2087	: Soma_AMA3_1 PORT MAP(
	A=> C(	2151	),
	B=>E(	1992	),
	Cin=> Carry( 	2086	),
	Cout=> Carry( 	2087	),
	S=> E(	2054	));
			
  U2088	: Soma_AMA3_1 PORT MAP(
	A=> C(	2152	),
	B=>E(	1993	),
	Cin=> Carry( 	2087	),
	Cout=> Carry( 	2088	),
	S=> E(	2055	));
			
  U2089	: Soma_AMA3_1 PORT MAP(
	A=> C(	2153	),
	B=>E(	1994	),
	Cin=> Carry( 	2088	),
	Cout=> Carry( 	2089	),
	S=> E(	2056	));
			
  U2090	: Soma_AMA3_1 PORT MAP(
	A=> C(	2154	),
	B=>E(	1995	),
	Cin=> Carry( 	2089	),
	Cout=> Carry( 	2090	),
	S=> E(	2057	));
			
  U2091	: Soma_AMA3_1 PORT MAP(
	A=> C(	2155	),
	B=>E(	1996	),
	Cin=> Carry( 	2090	),
	Cout=> Carry( 	2091	),
	S=> E(	2058	));
			
  U2092	: Soma_AMA3_1 PORT MAP(
	A=> C(	2156	),
	B=>E(	1997	),
	Cin=> Carry( 	2091	),
	Cout=> Carry( 	2092	),
	S=> E(	2059	));
			
  U2093	: Soma_AMA3_1 PORT MAP(
	A=> C(	2157	),
	B=>E(	1998	),
	Cin=> Carry( 	2092	),
	Cout=> Carry( 	2093	),
	S=> E(	2060	));
			
  U2094	: Soma_AMA3_1 PORT MAP(
	A=> C(	2158	),
	B=>E(	1999	),
	Cin=> Carry( 	2093	),
	Cout=> Carry( 	2094	),
	S=> E(	2061	));
			
  U2095	: Soma_AMA3_1 PORT MAP(
	A=> C(	2159	),
	B=>E(	2000	),
	Cin=> Carry( 	2094	),
	Cout=> Carry( 	2095	),
	S=> E(	2062	));
			
  U2096	: Soma_AMA3_1 PORT MAP(
	A=> C(	2160	),
	B=>E(	2001	),
	Cin=> Carry( 	2095	),
	Cout=> Carry( 	2096	),
	S=> E(	2063	));
			
  U2097	: Soma_AMA3_1 PORT MAP(
	A=> C(	2161	),
	B=>E(	2002	),
	Cin=> Carry( 	2096	),
	Cout=> Carry( 	2097	),
	S=> E(	2064	));
			
  U2098	: Soma_AMA3_1 PORT MAP(
	A=> C(	2162	),
	B=>E(	2003	),
	Cin=> Carry( 	2097	),
	Cout=> Carry( 	2098	),
	S=> E(	2065	));
			
  U2099	: Soma_AMA3_1 PORT MAP(
	A=> C(	2163	),
	B=>E(	2004	),
	Cin=> Carry( 	2098	),
	Cout=> Carry( 	2099	),
	S=> E(	2066	));
			
  U2100	: Soma_AMA3_1 PORT MAP(
	A=> C(	2164	),
	B=>E(	2005	),
	Cin=> Carry( 	2099	),
	Cout=> Carry( 	2100	),
	S=> E(	2067	));
			
  U2101	: Soma_AMA3_1 PORT MAP(
	A=> C(	2165	),
	B=>E(	2006	),
	Cin=> Carry( 	2100	),
	Cout=> Carry( 	2101	),
	S=> E(	2068	));
			
  U2102	: Soma_AMA3_1 PORT MAP(
	A=> C(	2166	),
	B=>E(	2007	),
	Cin=> Carry( 	2101	),
	Cout=> Carry( 	2102	),
	S=> E(	2069	));
			
  U2103	: Soma_AMA3_1 PORT MAP(
	A=> C(	2167	),
	B=>E(	2008	),
	Cin=> Carry( 	2102	),
	Cout=> Carry( 	2103	),
	S=> E(	2070	));
			
  U2104	: Soma_AMA3_1 PORT MAP(
	A=> C(	2168	),
	B=>E(	2009	),
	Cin=> Carry( 	2103	),
	Cout=> Carry( 	2104	),
	S=> E(	2071	));
			
  U2105	: Soma_AMA3_1 PORT MAP(
	A=> C(	2169	),
	B=>E(	2010	),
	Cin=> Carry( 	2104	),
	Cout=> Carry( 	2105	),
	S=> E(	2072	));
			
  U2106	: Soma_AMA3_1 PORT MAP(
	A=> C(	2170	),
	B=>E(	2011	),
	Cin=> Carry( 	2105	),
	Cout=> Carry( 	2106	),
	S=> E(	2073	));
			
  U2107	: Soma_AMA3_1 PORT MAP(
	A=> C(	2171	),
	B=>E(	2012	),
	Cin=> Carry( 	2106	),
	Cout=> Carry( 	2107	),
	S=> E(	2074	));
			
  U2108	: Soma_AMA3_1 PORT MAP(
	A=> C(	2172	),
	B=>E(	2013	),
	Cin=> Carry( 	2107	),
	Cout=> Carry( 	2108	),
	S=> E(	2075	));
			
  U2109	: Soma_AMA3_1 PORT MAP(
	A=> C(	2173	),
	B=>E(	2014	),
	Cin=> Carry( 	2108	),
	Cout=> Carry( 	2109	),
	S=> E(	2076	));
			
  U2110	: Soma_AMA3_1 PORT MAP(
	A=> C(	2174	),
	B=>E(	2015	),
	Cin=> Carry( 	2109	),
	Cout=> Carry( 	2110	),
	S=> E(	2077	));
			
  U2111	: Soma_AMA3_1 PORT MAP(
	A=> C(	2175	),
	B=>Carry(	2047	),
	Cin=> Carry( 	2110	),
	Cout=> Carry( 	2111	),
	S=> E(	2078	));

			
  U2112	: Soma_AMA3_1 PORT MAP(
	A=> C(	2176	),
	B=>E(	2016	),
	Cin=> '0'	,
	Cout=> Carry( 	2112	),
	S=> R(	34	));
			
  U2113	: Soma_AMA3_1 PORT MAP(
	A=> C(	2177	),
	B=>E(	2017	),
	Cin=> Carry( 	2112	),
	Cout=> Carry( 	2113	),
	S=> E(	2079	));
			
  U2114	: Soma_AMA3_1 PORT MAP(
	A=> C(	2178	),
	B=>E(	2018	),
	Cin=> Carry( 	2113	),
	Cout=> Carry( 	2114	),
	S=> E(	2080	));
			
  U2115	: Soma_AMA3_1 PORT MAP(
	A=> C(	2179	),
	B=>E(	2019	),
	Cin=> Carry( 	2114	),
	Cout=> Carry( 	2115	),
	S=> E(	2081	));
			
  U2116	: Soma_AMA3_1 PORT MAP(
	A=> C(	2180	),
	B=>E(	2020	),
	Cin=> Carry( 	2115	),
	Cout=> Carry( 	2116	),
	S=> E(	2082	));
			
  U2117	: Soma_AMA3_1 PORT MAP(
	A=> C(	2181	),
	B=>E(	2021	),
	Cin=> Carry( 	2116	),
	Cout=> Carry( 	2117	),
	S=> E(	2083	));
			
  U2118	: Soma_AMA3_1 PORT MAP(
	A=> C(	2182	),
	B=>E(	2022	),
	Cin=> Carry( 	2117	),
	Cout=> Carry( 	2118	),
	S=> E(	2084	));
			
  U2119	: Soma_AMA3_1 PORT MAP(
	A=> C(	2183	),
	B=>E(	2023	),
	Cin=> Carry( 	2118	),
	Cout=> Carry( 	2119	),
	S=> E(	2085	));
			
  U2120	: Soma_AMA3_1 PORT MAP(
	A=> C(	2184	),
	B=>E(	2024	),
	Cin=> Carry( 	2119	),
	Cout=> Carry( 	2120	),
	S=> E(	2086	));
			
  U2121	: Soma_AMA3_1 PORT MAP(
	A=> C(	2185	),
	B=>E(	2025	),
	Cin=> Carry( 	2120	),
	Cout=> Carry( 	2121	),
	S=> E(	2087	));
			
  U2122	: Soma_AMA3_1 PORT MAP(
	A=> C(	2186	),
	B=>E(	2026	),
	Cin=> Carry( 	2121	),
	Cout=> Carry( 	2122	),
	S=> E(	2088	));
			
  U2123	: Soma_AMA3_1 PORT MAP(
	A=> C(	2187	),
	B=>E(	2027	),
	Cin=> Carry( 	2122	),
	Cout=> Carry( 	2123	),
	S=> E(	2089	));
			
  U2124	: Soma_AMA3_1 PORT MAP(
	A=> C(	2188	),
	B=>E(	2028	),
	Cin=> Carry( 	2123	),
	Cout=> Carry( 	2124	),
	S=> E(	2090	));
			
  U2125	: Soma_AMA3_1 PORT MAP(
	A=> C(	2189	),
	B=>E(	2029	),
	Cin=> Carry( 	2124	),
	Cout=> Carry( 	2125	),
	S=> E(	2091	));
			
  U2126	: Soma_AMA3_1 PORT MAP(
	A=> C(	2190	),
	B=>E(	2030	),
	Cin=> Carry( 	2125	),
	Cout=> Carry( 	2126	),
	S=> E(	2092	));
			
  U2127	: Soma_AMA3_1 PORT MAP(
	A=> C(	2191	),
	B=>E(	2031	),
	Cin=> Carry( 	2126	),
	Cout=> Carry( 	2127	),
	S=> E(	2093	));
			
  U2128	: Soma_AMA3_1 PORT MAP(
	A=> C(	2192	),
	B=>E(	2032	),
	Cin=> Carry( 	2127	),
	Cout=> Carry( 	2128	),
	S=> E(	2094	));
			
  U2129	: Soma_AMA3_1 PORT MAP(
	A=> C(	2193	),
	B=>E(	2033	),
	Cin=> Carry( 	2128	),
	Cout=> Carry( 	2129	),
	S=> E(	2095	));
			
  U2130	: Soma_AMA3_1 PORT MAP(
	A=> C(	2194	),
	B=>E(	2034	),
	Cin=> Carry( 	2129	),
	Cout=> Carry( 	2130	),
	S=> E(	2096	));
			
  U2131	: Soma_AMA3_1 PORT MAP(
	A=> C(	2195	),
	B=>E(	2035	),
	Cin=> Carry( 	2130	),
	Cout=> Carry( 	2131	),
	S=> E(	2097	));
			
  U2132	: Soma_AMA3_1 PORT MAP(
	A=> C(	2196	),
	B=>E(	2036	),
	Cin=> Carry( 	2131	),
	Cout=> Carry( 	2132	),
	S=> E(	2098	));
			
  U2133	: Soma_AMA3_1 PORT MAP(
	A=> C(	2197	),
	B=>E(	2037	),
	Cin=> Carry( 	2132	),
	Cout=> Carry( 	2133	),
	S=> E(	2099	));
			
  U2134	: Soma_AMA3_1 PORT MAP(
	A=> C(	2198	),
	B=>E(	2038	),
	Cin=> Carry( 	2133	),
	Cout=> Carry( 	2134	),
	S=> E(	2100	));
			
  U2135	: Soma_AMA3_1 PORT MAP(
	A=> C(	2199	),
	B=>E(	2039	),
	Cin=> Carry( 	2134	),
	Cout=> Carry( 	2135	),
	S=> E(	2101	));
			
  U2136	: Soma_AMA3_1 PORT MAP(
	A=> C(	2200	),
	B=>E(	2040	),
	Cin=> Carry( 	2135	),
	Cout=> Carry( 	2136	),
	S=> E(	2102	));
			
  U2137	: Soma_AMA3_1 PORT MAP(
	A=> C(	2201	),
	B=>E(	2041	),
	Cin=> Carry( 	2136	),
	Cout=> Carry( 	2137	),
	S=> E(	2103	));
			
  U2138	: Soma_AMA3_1 PORT MAP(
	A=> C(	2202	),
	B=>E(	2042	),
	Cin=> Carry( 	2137	),
	Cout=> Carry( 	2138	),
	S=> E(	2104	));
			
  U2139	: Soma_AMA3_1 PORT MAP(
	A=> C(	2203	),
	B=>E(	2043	),
	Cin=> Carry( 	2138	),
	Cout=> Carry( 	2139	),
	S=> E(	2105	));
			
  U2140	: Soma_AMA3_1 PORT MAP(
	A=> C(	2204	),
	B=>E(	2044	),
	Cin=> Carry( 	2139	),
	Cout=> Carry( 	2140	),
	S=> E(	2106	));
			
  U2141	: Soma_AMA3_1 PORT MAP(
	A=> C(	2205	),
	B=>E(	2045	),
	Cin=> Carry( 	2140	),
	Cout=> Carry( 	2141	),
	S=> E(	2107	));
			
  U2142	: Soma_AMA3_1 PORT MAP(
	A=> C(	2206	),
	B=>E(	2046	),
	Cin=> Carry( 	2141	),
	Cout=> Carry( 	2142	),
	S=> E(	2108	));
			
  U2143	: Soma_AMA3_1 PORT MAP(
	A=> C(	2207	),
	B=>E(	2047	),
	Cin=> Carry( 	2142	),
	Cout=> Carry( 	2143	),
	S=> E(	2109	));
			
  U2144	: Soma_AMA3_1 PORT MAP(
	A=> C(	2208	),
	B=>E(	2048	),
	Cin=> Carry( 	2143	),
	Cout=> Carry( 	2144	),
	S=> E(	2110	));
			
  U2145	: Soma_AMA3_1 PORT MAP(
	A=> C(	2209	),
	B=>E(	2049	),
	Cin=> Carry( 	2144	),
	Cout=> Carry( 	2145	),
	S=> E(	2111	));
			
  U2146	: Soma_AMA3_1 PORT MAP(
	A=> C(	2210	),
	B=>E(	2050	),
	Cin=> Carry( 	2145	),
	Cout=> Carry( 	2146	),
	S=> E(	2112	));
			
  U2147	: Soma_AMA3_1 PORT MAP(
	A=> C(	2211	),
	B=>E(	2051	),
	Cin=> Carry( 	2146	),
	Cout=> Carry( 	2147	),
	S=> E(	2113	));
			
  U2148	: Soma_AMA3_1 PORT MAP(
	A=> C(	2212	),
	B=>E(	2052	),
	Cin=> Carry( 	2147	),
	Cout=> Carry( 	2148	),
	S=> E(	2114	));
			
  U2149	: Soma_AMA3_1 PORT MAP(
	A=> C(	2213	),
	B=>E(	2053	),
	Cin=> Carry( 	2148	),
	Cout=> Carry( 	2149	),
	S=> E(	2115	));
			
  U2150	: Soma_AMA3_1 PORT MAP(
	A=> C(	2214	),
	B=>E(	2054	),
	Cin=> Carry( 	2149	),
	Cout=> Carry( 	2150	),
	S=> E(	2116	));
			
  U2151	: Soma_AMA3_1 PORT MAP(
	A=> C(	2215	),
	B=>E(	2055	),
	Cin=> Carry( 	2150	),
	Cout=> Carry( 	2151	),
	S=> E(	2117	));
			
  U2152	: Soma_AMA3_1 PORT MAP(
	A=> C(	2216	),
	B=>E(	2056	),
	Cin=> Carry( 	2151	),
	Cout=> Carry( 	2152	),
	S=> E(	2118	));
			
  U2153	: Soma_AMA3_1 PORT MAP(
	A=> C(	2217	),
	B=>E(	2057	),
	Cin=> Carry( 	2152	),
	Cout=> Carry( 	2153	),
	S=> E(	2119	));
			
  U2154	: Soma_AMA3_1 PORT MAP(
	A=> C(	2218	),
	B=>E(	2058	),
	Cin=> Carry( 	2153	),
	Cout=> Carry( 	2154	),
	S=> E(	2120	));
			
  U2155	: Soma_AMA3_1 PORT MAP(
	A=> C(	2219	),
	B=>E(	2059	),
	Cin=> Carry( 	2154	),
	Cout=> Carry( 	2155	),
	S=> E(	2121	));
			
  U2156	: Soma_AMA3_1 PORT MAP(
	A=> C(	2220	),
	B=>E(	2060	),
	Cin=> Carry( 	2155	),
	Cout=> Carry( 	2156	),
	S=> E(	2122	));
			
  U2157	: Soma_AMA3_1 PORT MAP(
	A=> C(	2221	),
	B=>E(	2061	),
	Cin=> Carry( 	2156	),
	Cout=> Carry( 	2157	),
	S=> E(	2123	));
			
  U2158	: Soma_AMA3_1 PORT MAP(
	A=> C(	2222	),
	B=>E(	2062	),
	Cin=> Carry( 	2157	),
	Cout=> Carry( 	2158	),
	S=> E(	2124	));
			
  U2159	: Soma_AMA3_1 PORT MAP(
	A=> C(	2223	),
	B=>E(	2063	),
	Cin=> Carry( 	2158	),
	Cout=> Carry( 	2159	),
	S=> E(	2125	));
			
  U2160	: Soma_AMA3_1 PORT MAP(
	A=> C(	2224	),
	B=>E(	2064	),
	Cin=> Carry( 	2159	),
	Cout=> Carry( 	2160	),
	S=> E(	2126	));
			
  U2161	: Soma_AMA3_1 PORT MAP(
	A=> C(	2225	),
	B=>E(	2065	),
	Cin=> Carry( 	2160	),
	Cout=> Carry( 	2161	),
	S=> E(	2127	));
			
  U2162	: Soma_AMA3_1 PORT MAP(
	A=> C(	2226	),
	B=>E(	2066	),
	Cin=> Carry( 	2161	),
	Cout=> Carry( 	2162	),
	S=> E(	2128	));
			
  U2163	: Soma_AMA3_1 PORT MAP(
	A=> C(	2227	),
	B=>E(	2067	),
	Cin=> Carry( 	2162	),
	Cout=> Carry( 	2163	),
	S=> E(	2129	));
			
  U2164	: Soma_AMA3_1 PORT MAP(
	A=> C(	2228	),
	B=>E(	2068	),
	Cin=> Carry( 	2163	),
	Cout=> Carry( 	2164	),
	S=> E(	2130	));
			
  U2165	: Soma_AMA3_1 PORT MAP(
	A=> C(	2229	),
	B=>E(	2069	),
	Cin=> Carry( 	2164	),
	Cout=> Carry( 	2165	),
	S=> E(	2131	));
			
  U2166	: Soma_AMA3_1 PORT MAP(
	A=> C(	2230	),
	B=>E(	2070	),
	Cin=> Carry( 	2165	),
	Cout=> Carry( 	2166	),
	S=> E(	2132	));
			
  U2167	: Soma_AMA3_1 PORT MAP(
	A=> C(	2231	),
	B=>E(	2071	),
	Cin=> Carry( 	2166	),
	Cout=> Carry( 	2167	),
	S=> E(	2133	));
			
  U2168	: Soma_AMA3_1 PORT MAP(
	A=> C(	2232	),
	B=>E(	2072	),
	Cin=> Carry( 	2167	),
	Cout=> Carry( 	2168	),
	S=> E(	2134	));
			
  U2169	: Soma_AMA3_1 PORT MAP(
	A=> C(	2233	),
	B=>E(	2073	),
	Cin=> Carry( 	2168	),
	Cout=> Carry( 	2169	),
	S=> E(	2135	));
			
  U2170	: Soma_AMA3_1 PORT MAP(
	A=> C(	2234	),
	B=>E(	2074	),
	Cin=> Carry( 	2169	),
	Cout=> Carry( 	2170	),
	S=> E(	2136	));
			
  U2171	: Soma_AMA3_1 PORT MAP(
	A=> C(	2235	),
	B=>E(	2075	),
	Cin=> Carry( 	2170	),
	Cout=> Carry( 	2171	),
	S=> E(	2137	));
			
  U2172	: Soma_AMA3_1 PORT MAP(
	A=> C(	2236	),
	B=>E(	2076	),
	Cin=> Carry( 	2171	),
	Cout=> Carry( 	2172	),
	S=> E(	2138	));
			
  U2173	: Soma_AMA3_1 PORT MAP(
	A=> C(	2237	),
	B=>E(	2077	),
	Cin=> Carry( 	2172	),
	Cout=> Carry( 	2173	),
	S=> E(	2139	));
			
  U2174	: Soma_AMA3_1 PORT MAP(
	A=> C(	2238	),
	B=>E(	2078	),
	Cin=> Carry( 	2173	),
	Cout=> Carry( 	2174	),
	S=> E(	2140	));
			
  U2175	: Soma_AMA3_1 PORT MAP(
	A=> C(	2239	),
	B=>Carry(	2111	),
	Cin=> Carry( 	2174	),
	Cout=> Carry( 	2175	),
	S=> E(	2141	));

			
  U2176	: Soma_AMA3_1 PORT MAP(
	A=> C(	2240	),
	B=>E(	2079	),
	Cin=> '0'	,
	Cout=> Carry( 	2176	),
	S=> R(	35	));
			
  U2177	: Soma_AMA3_1 PORT MAP(
	A=> C(	2241	),
	B=>E(	2080	),
	Cin=> Carry( 	2176	),
	Cout=> Carry( 	2177	),
	S=> E(	2142	));
			
  U2178	: Soma_AMA3_1 PORT MAP(
	A=> C(	2242	),
	B=>E(	2081	),
	Cin=> Carry( 	2177	),
	Cout=> Carry( 	2178	),
	S=> E(	2143	));
			
  U2179	: Soma_AMA3_1 PORT MAP(
	A=> C(	2243	),
	B=>E(	2082	),
	Cin=> Carry( 	2178	),
	Cout=> Carry( 	2179	),
	S=> E(	2144	));
			
  U2180	: Soma_AMA3_1 PORT MAP(
	A=> C(	2244	),
	B=>E(	2083	),
	Cin=> Carry( 	2179	),
	Cout=> Carry( 	2180	),
	S=> E(	2145	));
			
  U2181	: Soma_AMA3_1 PORT MAP(
	A=> C(	2245	),
	B=>E(	2084	),
	Cin=> Carry( 	2180	),
	Cout=> Carry( 	2181	),
	S=> E(	2146	));
			
  U2182	: Soma_AMA3_1 PORT MAP(
	A=> C(	2246	),
	B=>E(	2085	),
	Cin=> Carry( 	2181	),
	Cout=> Carry( 	2182	),
	S=> E(	2147	));
			
  U2183	: Soma_AMA3_1 PORT MAP(
	A=> C(	2247	),
	B=>E(	2086	),
	Cin=> Carry( 	2182	),
	Cout=> Carry( 	2183	),
	S=> E(	2148	));
			
  U2184	: Soma_AMA3_1 PORT MAP(
	A=> C(	2248	),
	B=>E(	2087	),
	Cin=> Carry( 	2183	),
	Cout=> Carry( 	2184	),
	S=> E(	2149	));
			
  U2185	: Soma_AMA3_1 PORT MAP(
	A=> C(	2249	),
	B=>E(	2088	),
	Cin=> Carry( 	2184	),
	Cout=> Carry( 	2185	),
	S=> E(	2150	));
			
  U2186	: Soma_AMA3_1 PORT MAP(
	A=> C(	2250	),
	B=>E(	2089	),
	Cin=> Carry( 	2185	),
	Cout=> Carry( 	2186	),
	S=> E(	2151	));
			
  U2187	: Soma_AMA3_1 PORT MAP(
	A=> C(	2251	),
	B=>E(	2090	),
	Cin=> Carry( 	2186	),
	Cout=> Carry( 	2187	),
	S=> E(	2152	));
			
  U2188	: Soma_AMA3_1 PORT MAP(
	A=> C(	2252	),
	B=>E(	2091	),
	Cin=> Carry( 	2187	),
	Cout=> Carry( 	2188	),
	S=> E(	2153	));
			
  U2189	: Soma_AMA3_1 PORT MAP(
	A=> C(	2253	),
	B=>E(	2092	),
	Cin=> Carry( 	2188	),
	Cout=> Carry( 	2189	),
	S=> E(	2154	));
			
  U2190	: Soma_AMA3_1 PORT MAP(
	A=> C(	2254	),
	B=>E(	2093	),
	Cin=> Carry( 	2189	),
	Cout=> Carry( 	2190	),
	S=> E(	2155	));
			
  U2191	: Soma_AMA3_1 PORT MAP(
	A=> C(	2255	),
	B=>E(	2094	),
	Cin=> Carry( 	2190	),
	Cout=> Carry( 	2191	),
	S=> E(	2156	));
			
  U2192	: Soma_AMA3_1 PORT MAP(
	A=> C(	2256	),
	B=>E(	2095	),
	Cin=> Carry( 	2191	),
	Cout=> Carry( 	2192	),
	S=> E(	2157	));
			
  U2193	: Soma_AMA3_1 PORT MAP(
	A=> C(	2257	),
	B=>E(	2096	),
	Cin=> Carry( 	2192	),
	Cout=> Carry( 	2193	),
	S=> E(	2158	));
			
  U2194	: Soma_AMA3_1 PORT MAP(
	A=> C(	2258	),
	B=>E(	2097	),
	Cin=> Carry( 	2193	),
	Cout=> Carry( 	2194	),
	S=> E(	2159	));
			
  U2195	: Soma_AMA3_1 PORT MAP(
	A=> C(	2259	),
	B=>E(	2098	),
	Cin=> Carry( 	2194	),
	Cout=> Carry( 	2195	),
	S=> E(	2160	));
			
  U2196	: Soma_AMA3_1 PORT MAP(
	A=> C(	2260	),
	B=>E(	2099	),
	Cin=> Carry( 	2195	),
	Cout=> Carry( 	2196	),
	S=> E(	2161	));
			
  U2197	: Soma_AMA3_1 PORT MAP(
	A=> C(	2261	),
	B=>E(	2100	),
	Cin=> Carry( 	2196	),
	Cout=> Carry( 	2197	),
	S=> E(	2162	));
			
  U2198	: Soma_AMA3_1 PORT MAP(
	A=> C(	2262	),
	B=>E(	2101	),
	Cin=> Carry( 	2197	),
	Cout=> Carry( 	2198	),
	S=> E(	2163	));
			
  U2199	: Soma_AMA3_1 PORT MAP(
	A=> C(	2263	),
	B=>E(	2102	),
	Cin=> Carry( 	2198	),
	Cout=> Carry( 	2199	),
	S=> E(	2164	));
			
  U2200	: Soma_AMA3_1 PORT MAP(
	A=> C(	2264	),
	B=>E(	2103	),
	Cin=> Carry( 	2199	),
	Cout=> Carry( 	2200	),
	S=> E(	2165	));
			
  U2201	: Soma_AMA3_1 PORT MAP(
	A=> C(	2265	),
	B=>E(	2104	),
	Cin=> Carry( 	2200	),
	Cout=> Carry( 	2201	),
	S=> E(	2166	));
			
  U2202	: Soma_AMA3_1 PORT MAP(
	A=> C(	2266	),
	B=>E(	2105	),
	Cin=> Carry( 	2201	),
	Cout=> Carry( 	2202	),
	S=> E(	2167	));
			
  U2203	: Soma_AMA3_1 PORT MAP(
	A=> C(	2267	),
	B=>E(	2106	),
	Cin=> Carry( 	2202	),
	Cout=> Carry( 	2203	),
	S=> E(	2168	));
			
  U2204	: Soma_AMA3_1 PORT MAP(
	A=> C(	2268	),
	B=>E(	2107	),
	Cin=> Carry( 	2203	),
	Cout=> Carry( 	2204	),
	S=> E(	2169	));
			
  U2205	: Soma_AMA3_1 PORT MAP(
	A=> C(	2269	),
	B=>E(	2108	),
	Cin=> Carry( 	2204	),
	Cout=> Carry( 	2205	),
	S=> E(	2170	));
			
  U2206	: Soma_AMA3_1 PORT MAP(
	A=> C(	2270	),
	B=>E(	2109	),
	Cin=> Carry( 	2205	),
	Cout=> Carry( 	2206	),
	S=> E(	2171	));
			
  U2207	: Soma_AMA3_1 PORT MAP(
	A=> C(	2271	),
	B=>E(	2110	),
	Cin=> Carry( 	2206	),
	Cout=> Carry( 	2207	),
	S=> E(	2172	));
			
  U2208	: Soma_AMA3_1 PORT MAP(
	A=> C(	2272	),
	B=>E(	2111	),
	Cin=> Carry( 	2207	),
	Cout=> Carry( 	2208	),
	S=> E(	2173	));
			
  U2209	: Soma_AMA3_1 PORT MAP(
	A=> C(	2273	),
	B=>E(	2112	),
	Cin=> Carry( 	2208	),
	Cout=> Carry( 	2209	),
	S=> E(	2174	));
			
  U2210	: Soma_AMA3_1 PORT MAP(
	A=> C(	2274	),
	B=>E(	2113	),
	Cin=> Carry( 	2209	),
	Cout=> Carry( 	2210	),
	S=> E(	2175	));
			
  U2211	: Soma_AMA3_1 PORT MAP(
	A=> C(	2275	),
	B=>E(	2114	),
	Cin=> Carry( 	2210	),
	Cout=> Carry( 	2211	),
	S=> E(	2176	));
			
  U2212	: Soma_AMA3_1 PORT MAP(
	A=> C(	2276	),
	B=>E(	2115	),
	Cin=> Carry( 	2211	),
	Cout=> Carry( 	2212	),
	S=> E(	2177	));
			
  U2213	: Soma_AMA3_1 PORT MAP(
	A=> C(	2277	),
	B=>E(	2116	),
	Cin=> Carry( 	2212	),
	Cout=> Carry( 	2213	),
	S=> E(	2178	));
			
  U2214	: Soma_AMA3_1 PORT MAP(
	A=> C(	2278	),
	B=>E(	2117	),
	Cin=> Carry( 	2213	),
	Cout=> Carry( 	2214	),
	S=> E(	2179	));
			
  U2215	: Soma_AMA3_1 PORT MAP(
	A=> C(	2279	),
	B=>E(	2118	),
	Cin=> Carry( 	2214	),
	Cout=> Carry( 	2215	),
	S=> E(	2180	));
			
  U2216	: Soma_AMA3_1 PORT MAP(
	A=> C(	2280	),
	B=>E(	2119	),
	Cin=> Carry( 	2215	),
	Cout=> Carry( 	2216	),
	S=> E(	2181	));
			
  U2217	: Soma_AMA3_1 PORT MAP(
	A=> C(	2281	),
	B=>E(	2120	),
	Cin=> Carry( 	2216	),
	Cout=> Carry( 	2217	),
	S=> E(	2182	));
			
  U2218	: Soma_AMA3_1 PORT MAP(
	A=> C(	2282	),
	B=>E(	2121	),
	Cin=> Carry( 	2217	),
	Cout=> Carry( 	2218	),
	S=> E(	2183	));
			
  U2219	: Soma_AMA3_1 PORT MAP(
	A=> C(	2283	),
	B=>E(	2122	),
	Cin=> Carry( 	2218	),
	Cout=> Carry( 	2219	),
	S=> E(	2184	));
			
  U2220	: Soma_AMA3_1 PORT MAP(
	A=> C(	2284	),
	B=>E(	2123	),
	Cin=> Carry( 	2219	),
	Cout=> Carry( 	2220	),
	S=> E(	2185	));
			
  U2221	: Soma_AMA3_1 PORT MAP(
	A=> C(	2285	),
	B=>E(	2124	),
	Cin=> Carry( 	2220	),
	Cout=> Carry( 	2221	),
	S=> E(	2186	));
			
  U2222	: Soma_AMA3_1 PORT MAP(
	A=> C(	2286	),
	B=>E(	2125	),
	Cin=> Carry( 	2221	),
	Cout=> Carry( 	2222	),
	S=> E(	2187	));
			
  U2223	: Soma_AMA3_1 PORT MAP(
	A=> C(	2287	),
	B=>E(	2126	),
	Cin=> Carry( 	2222	),
	Cout=> Carry( 	2223	),
	S=> E(	2188	));
			
  U2224	: Soma_AMA3_1 PORT MAP(
	A=> C(	2288	),
	B=>E(	2127	),
	Cin=> Carry( 	2223	),
	Cout=> Carry( 	2224	),
	S=> E(	2189	));
			
  U2225	: Soma_AMA3_1 PORT MAP(
	A=> C(	2289	),
	B=>E(	2128	),
	Cin=> Carry( 	2224	),
	Cout=> Carry( 	2225	),
	S=> E(	2190	));
			
  U2226	: Soma_AMA3_1 PORT MAP(
	A=> C(	2290	),
	B=>E(	2129	),
	Cin=> Carry( 	2225	),
	Cout=> Carry( 	2226	),
	S=> E(	2191	));
			
  U2227	: Soma_AMA3_1 PORT MAP(
	A=> C(	2291	),
	B=>E(	2130	),
	Cin=> Carry( 	2226	),
	Cout=> Carry( 	2227	),
	S=> E(	2192	));
			
  U2228	: Soma_AMA3_1 PORT MAP(
	A=> C(	2292	),
	B=>E(	2131	),
	Cin=> Carry( 	2227	),
	Cout=> Carry( 	2228	),
	S=> E(	2193	));
			
  U2229	: Soma_AMA3_1 PORT MAP(
	A=> C(	2293	),
	B=>E(	2132	),
	Cin=> Carry( 	2228	),
	Cout=> Carry( 	2229	),
	S=> E(	2194	));
			
  U2230	: Soma_AMA3_1 PORT MAP(
	A=> C(	2294	),
	B=>E(	2133	),
	Cin=> Carry( 	2229	),
	Cout=> Carry( 	2230	),
	S=> E(	2195	));
			
  U2231	: Soma_AMA3_1 PORT MAP(
	A=> C(	2295	),
	B=>E(	2134	),
	Cin=> Carry( 	2230	),
	Cout=> Carry( 	2231	),
	S=> E(	2196	));
			
  U2232	: Soma_AMA3_1 PORT MAP(
	A=> C(	2296	),
	B=>E(	2135	),
	Cin=> Carry( 	2231	),
	Cout=> Carry( 	2232	),
	S=> E(	2197	));
			
  U2233	: Soma_AMA3_1 PORT MAP(
	A=> C(	2297	),
	B=>E(	2136	),
	Cin=> Carry( 	2232	),
	Cout=> Carry( 	2233	),
	S=> E(	2198	));
			
  U2234	: Soma_AMA3_1 PORT MAP(
	A=> C(	2298	),
	B=>E(	2137	),
	Cin=> Carry( 	2233	),
	Cout=> Carry( 	2234	),
	S=> E(	2199	));
			
  U2235	: Soma_AMA3_1 PORT MAP(
	A=> C(	2299	),
	B=>E(	2138	),
	Cin=> Carry( 	2234	),
	Cout=> Carry( 	2235	),
	S=> E(	2200	));
			
  U2236	: Soma_AMA3_1 PORT MAP(
	A=> C(	2300	),
	B=>E(	2139	),
	Cin=> Carry( 	2235	),
	Cout=> Carry( 	2236	),
	S=> E(	2201	));
			
  U2237	: Soma_AMA3_1 PORT MAP(
	A=> C(	2301	),
	B=>E(	2140	),
	Cin=> Carry( 	2236	),
	Cout=> Carry( 	2237	),
	S=> E(	2202	));
			
  U2238	: Soma_AMA3_1 PORT MAP(
	A=> C(	2302	),
	B=>E(	2141	),
	Cin=> Carry( 	2237	),
	Cout=> Carry( 	2238	),
	S=> E(	2203	));
			
  U2239	: Soma_AMA3_1 PORT MAP(
	A=> C(	2303	),
	B=>Carry(	2175	),
	Cin=> Carry( 	2238	),
	Cout=> Carry( 	2239	),
	S=> E(	2204	));

			
  U2240	: Soma_AMA3_1 PORT MAP(
	A=> C(	2304	),
	B=>E(	2142	),
	Cin=> '0'	,
	Cout=> Carry( 	2240	),
	S=> R(	36	));
			
  U2241	: Soma_AMA3_1 PORT MAP(
	A=> C(	2305	),
	B=>E(	2143	),
	Cin=> Carry( 	2240	),
	Cout=> Carry( 	2241	),
	S=> E(	2205	));
			
  U2242	: Soma_AMA3_1 PORT MAP(
	A=> C(	2306	),
	B=>E(	2144	),
	Cin=> Carry( 	2241	),
	Cout=> Carry( 	2242	),
	S=> E(	2206	));
			
  U2243	: Soma_AMA3_1 PORT MAP(
	A=> C(	2307	),
	B=>E(	2145	),
	Cin=> Carry( 	2242	),
	Cout=> Carry( 	2243	),
	S=> E(	2207	));
			
  U2244	: Soma_AMA3_1 PORT MAP(
	A=> C(	2308	),
	B=>E(	2146	),
	Cin=> Carry( 	2243	),
	Cout=> Carry( 	2244	),
	S=> E(	2208	));
			
  U2245	: Soma_AMA3_1 PORT MAP(
	A=> C(	2309	),
	B=>E(	2147	),
	Cin=> Carry( 	2244	),
	Cout=> Carry( 	2245	),
	S=> E(	2209	));
			
  U2246	: Soma_AMA3_1 PORT MAP(
	A=> C(	2310	),
	B=>E(	2148	),
	Cin=> Carry( 	2245	),
	Cout=> Carry( 	2246	),
	S=> E(	2210	));
			
  U2247	: Soma_AMA3_1 PORT MAP(
	A=> C(	2311	),
	B=>E(	2149	),
	Cin=> Carry( 	2246	),
	Cout=> Carry( 	2247	),
	S=> E(	2211	));
			
  U2248	: Soma_AMA3_1 PORT MAP(
	A=> C(	2312	),
	B=>E(	2150	),
	Cin=> Carry( 	2247	),
	Cout=> Carry( 	2248	),
	S=> E(	2212	));
			
  U2249	: Soma_AMA3_1 PORT MAP(
	A=> C(	2313	),
	B=>E(	2151	),
	Cin=> Carry( 	2248	),
	Cout=> Carry( 	2249	),
	S=> E(	2213	));
			
  U2250	: Soma_AMA3_1 PORT MAP(
	A=> C(	2314	),
	B=>E(	2152	),
	Cin=> Carry( 	2249	),
	Cout=> Carry( 	2250	),
	S=> E(	2214	));
			
  U2251	: Soma_AMA3_1 PORT MAP(
	A=> C(	2315	),
	B=>E(	2153	),
	Cin=> Carry( 	2250	),
	Cout=> Carry( 	2251	),
	S=> E(	2215	));
			
  U2252	: Soma_AMA3_1 PORT MAP(
	A=> C(	2316	),
	B=>E(	2154	),
	Cin=> Carry( 	2251	),
	Cout=> Carry( 	2252	),
	S=> E(	2216	));
			
  U2253	: Soma_AMA3_1 PORT MAP(
	A=> C(	2317	),
	B=>E(	2155	),
	Cin=> Carry( 	2252	),
	Cout=> Carry( 	2253	),
	S=> E(	2217	));
	
  U2254	: Soma_AMA3_1 PORT MAP(
	A=> C(	2318	),
	B=>E(	2156	),
	Cin=> Carry( 	2253	),
	Cout=> Carry( 	2254	),
	S=> E(	2218	));
			
  U2255	: Soma_AMA3_1 PORT MAP(
	A=> C(	2319	),
	B=>E(	2157	),
	Cin=> Carry( 	2254	),
	Cout=> Carry( 	2255	),
	S=> E(	2219	));
			
  U2256	: Soma_AMA3_1 PORT MAP(
	A=> C(	2320	),
	B=>E(	2158	),
	Cin=> Carry( 	2255	),
	Cout=> Carry( 	2256	),
	S=> E(	2220	));
			
  U2257	: Soma_AMA3_1 PORT MAP(
	A=> C(	2321	),
	B=>E(	2159	),
	Cin=> Carry( 	2256	),
	Cout=> Carry( 	2257	),
	S=> E(	2221	));
			
  U2258	: Soma_AMA3_1 PORT MAP(
	A=> C(	2322	),
	B=>E(	2160	),
	Cin=> Carry( 	2257	),
	Cout=> Carry( 	2258	),
	S=> E(	2222	));
			
  U2259	: Soma_AMA3_1 PORT MAP(
	A=> C(	2323	),
	B=>E(	2161	),
	Cin=> Carry( 	2258	),
	Cout=> Carry( 	2259	),
	S=> E(	2223	));
			
  U2260	: Soma_AMA3_1 PORT MAP(
	A=> C(	2324	),
	B=>E(	2162	),
	Cin=> Carry( 	2259	),
	Cout=> Carry( 	2260	),
	S=> E(	2224	));
			
  U2261	: Soma_AMA3_1 PORT MAP(
	A=> C(	2325	),
	B=>E(	2163	),
	Cin=> Carry( 	2260	),
	Cout=> Carry( 	2261	),
	S=> E(	2225	));
			
  U2262	: Soma_AMA3_1 PORT MAP(
	A=> C(	2326	),
	B=>E(	2164	),
	Cin=> Carry( 	2261	),
	Cout=> Carry( 	2262	),
	S=> E(	2226	));
			
  U2263	: Soma_AMA3_1 PORT MAP(
	A=> C(	2327	),
	B=>E(	2165	),
	Cin=> Carry( 	2262	),
	Cout=> Carry( 	2263	),
	S=> E(	2227	));
			
  U2264	: Soma_AMA3_1 PORT MAP(
	A=> C(	2328	),
	B=>E(	2166	),
	Cin=> Carry( 	2263	),
	Cout=> Carry( 	2264	),
	S=> E(	2228	));
			
  U2265	: Soma_AMA3_1 PORT MAP(
	A=> C(	2329	),
	B=>E(	2167	),
	Cin=> Carry( 	2264	),
	Cout=> Carry( 	2265	),
	S=> E(	2229	));
			
  U2266	: Soma_AMA3_1 PORT MAP(
	A=> C(	2330	),
	B=>E(	2168	),
	Cin=> Carry( 	2265	),
	Cout=> Carry( 	2266	),
	S=> E(	2230	));
			
  U2267	: Soma_AMA3_1 PORT MAP(
	A=> C(	2331	),
	B=>E(	2169	),
	Cin=> Carry( 	2266	),
	Cout=> Carry( 	2267	),
	S=> E(	2231	));
			
  U2268	: Soma_AMA3_1 PORT MAP(
	A=> C(	2332	),
	B=>E(	2170	),
	Cin=> Carry( 	2267	),
	Cout=> Carry( 	2268	),
	S=> E(	2232	));
			
  U2269	: Soma_AMA3_1 PORT MAP(
	A=> C(	2333	),
	B=>E(	2171	),
	Cin=> Carry( 	2268	),
	Cout=> Carry( 	2269	),
	S=> E(	2233	));
			
  U2270	: Soma_AMA3_1 PORT MAP(
	A=> C(	2334	),
	B=>E(	2172	),
	Cin=> Carry( 	2269	),
	Cout=> Carry( 	2270	),
	S=> E(	2234	));
			
  U2271	: Soma_AMA3_1 PORT MAP(
	A=> C(	2335	),
	B=>E(	2173	),
	Cin=> Carry( 	2270	),
	Cout=> Carry( 	2271	),
	S=> E(	2235	));
			
  U2272	: Soma_AMA3_1 PORT MAP(
	A=> C(	2336	),
	B=>E(	2174	),
	Cin=> Carry( 	2271	),
	Cout=> Carry( 	2272	),
	S=> E(	2236	));
			
  U2273	: Soma_AMA3_1 PORT MAP(
	A=> C(	2337	),
	B=>E(	2175	),
	Cin=> Carry( 	2272	),
	Cout=> Carry( 	2273	),
	S=> E(	2237	));
			
  U2274	: Soma_AMA3_1 PORT MAP(
	A=> C(	2338	),
	B=>E(	2176	),
	Cin=> Carry( 	2273	),
	Cout=> Carry( 	2274	),
	S=> E(	2238	));
			
  U2275	: Soma_AMA3_1 PORT MAP(
	A=> C(	2339	),
	B=>E(	2177	),
	Cin=> Carry( 	2274	),
	Cout=> Carry( 	2275	),
	S=> E(	2239	));
			
  U2276	: Soma_AMA3_1 PORT MAP(
	A=> C(	2340	),
	B=>E(	2178	),
	Cin=> Carry( 	2275	),
	Cout=> Carry( 	2276	),
	S=> E(	2240	));
			
  U2277	: Soma_AMA3_1 PORT MAP(
	A=> C(	2341	),
	B=>E(	2179	),
	Cin=> Carry( 	2276	),
	Cout=> Carry( 	2277	),
	S=> E(	2241	));
			
  U2278	: Soma_AMA3_1 PORT MAP(
	A=> C(	2342	),
	B=>E(	2180	),
	Cin=> Carry( 	2277	),
	Cout=> Carry( 	2278	),
	S=> E(	2242	));
			
  U2279	: Soma_AMA3_1 PORT MAP(
	A=> C(	2343	),
	B=>E(	2181	),
	Cin=> Carry( 	2278	),
	Cout=> Carry( 	2279	),
	S=> E(	2243	));
			
  U2280	: Soma_AMA3_1 PORT MAP(
	A=> C(	2344	),
	B=>E(	2182	),
	Cin=> Carry( 	2279	),
	Cout=> Carry( 	2280	),
	S=> E(	2244	));
			
  U2281	: Soma_AMA3_1 PORT MAP(
	A=> C(	2345	),
	B=>E(	2183	),
	Cin=> Carry( 	2280	),
	Cout=> Carry( 	2281	),
	S=> E(	2245	));
			
  U2282	: Soma_AMA3_1 PORT MAP(
	A=> C(	2346	),
	B=>E(	2184	),
	Cin=> Carry( 	2281	),
	Cout=> Carry( 	2282	),
	S=> E(	2246	));
			
  U2283	: Soma_AMA3_1 PORT MAP(
	A=> C(	2347	),
	B=>E(	2185	),
	Cin=> Carry( 	2282	),
	Cout=> Carry( 	2283	),
	S=> E(	2247	));
			
  U2284	: Soma_AMA3_1 PORT MAP(
	A=> C(	2348	),
	B=>E(	2186	),
	Cin=> Carry( 	2283	),
	Cout=> Carry( 	2284	),
	S=> E(	2248	));
			
  U2285	: Soma_AMA3_1 PORT MAP(
	A=> C(	2349	),
	B=>E(	2187	),
	Cin=> Carry( 	2284	),
	Cout=> Carry( 	2285	),
	S=> E(	2249	));
			
  U2286	: Soma_AMA3_1 PORT MAP(
	A=> C(	2350	),
	B=>E(	2188	),
	Cin=> Carry( 	2285	),
	Cout=> Carry( 	2286	),
	S=> E(	2250	));
			
  U2287	: Soma_AMA3_1 PORT MAP(
	A=> C(	2351	),
	B=>E(	2189	),
	Cin=> Carry( 	2286	),
	Cout=> Carry( 	2287	),
	S=> E(	2251	));
			
  U2288	: Soma_AMA3_1 PORT MAP(
	A=> C(	2352	),
	B=>E(	2190	),
	Cin=> Carry( 	2287	),
	Cout=> Carry( 	2288	),
	S=> E(	2252	));
			
  U2289	: Soma_AMA3_1 PORT MAP(
	A=> C(	2353	),
	B=>E(	2191	),
	Cin=> Carry( 	2288	),
	Cout=> Carry( 	2289	),
	S=> E(	2253	));
			
  U2290	: Soma_AMA3_1 PORT MAP(
	A=> C(	2354	),
	B=>E(	2192	),
	Cin=> Carry( 	2289	),
	Cout=> Carry( 	2290	),
	S=> E(	2254	));
			
  U2291	: Soma_AMA3_1 PORT MAP(
	A=> C(	2355	),
	B=>E(	2193	),
	Cin=> Carry( 	2290	),
	Cout=> Carry( 	2291	),
	S=> E(	2255	));
			
  U2292	: Soma_AMA3_1 PORT MAP(
	A=> C(	2356	),
	B=>E(	2194	),
	Cin=> Carry( 	2291	),
	Cout=> Carry( 	2292	),
	S=> E(	2256	));
			
  U2293	: Soma_AMA3_1 PORT MAP(
	A=> C(	2357	),
	B=>E(	2195	),
	Cin=> Carry( 	2292	),
	Cout=> Carry( 	2293	),
	S=> E(	2257	));
			
  U2294	: Soma_AMA3_1 PORT MAP(
	A=> C(	2358	),
	B=>E(	2196	),
	Cin=> Carry( 	2293	),
	Cout=> Carry( 	2294	),
	S=> E(	2258	));
			
  U2295	: Soma_AMA3_1 PORT MAP(
	A=> C(	2359	),
	B=>E(	2197	),
	Cin=> Carry( 	2294	),
	Cout=> Carry( 	2295	),
	S=> E(	2259	));
			
  U2296	: Soma_AMA3_1 PORT MAP(
	A=> C(	2360	),
	B=>E(	2198	),
	Cin=> Carry( 	2295	),
	Cout=> Carry( 	2296	),
	S=> E(	2260	));
			
  U2297	: Soma_AMA3_1 PORT MAP(
	A=> C(	2361	),
	B=>E(	2199	),
	Cin=> Carry( 	2296	),
	Cout=> Carry( 	2297	),
	S=> E(	2261	));
			
  U2298	: Soma_AMA3_1 PORT MAP(
	A=> C(	2362	),
	B=>E(	2200	),
	Cin=> Carry( 	2297	),
	Cout=> Carry( 	2298	),
	S=> E(	2262	));
			
  U2299	: Soma_AMA3_1 PORT MAP(
	A=> C(	2363	),
	B=>E(	2201	),
	Cin=> Carry( 	2298	),
	Cout=> Carry( 	2299	),
	S=> E(	2263	));
			
  U2300	: Soma_AMA3_1 PORT MAP(
	A=> C(	2364	),
	B=>E(	2202	),
	Cin=> Carry( 	2299	),
	Cout=> Carry( 	2300	),
	S=> E(	2264	));
			
  U2301	: Soma_AMA3_1 PORT MAP(
	A=> C(	2365	),
	B=>E(	2203	),
	Cin=> Carry( 	2300	),
	Cout=> Carry( 	2301	),
	S=> E(	2265	));
			
  U2302	: Soma_AMA3_1 PORT MAP(
	A=> C(	2366	),
	B=>E(	2204	),
	Cin=> Carry( 	2301	),
	Cout=> Carry( 	2302	),
	S=> E(	2266	));
			
  U2303	: Soma_AMA3_1 PORT MAP(
	A=> C(	2367	),
	B=>Carry(	2239	),
	Cin=> Carry( 	2302	),
	Cout=> Carry( 	2303	),
	S=> E(	2267	));

			
  U2304	: Soma_AMA3_1 PORT MAP(
	A=> C(	2368	),
	B=>E(	2205	),
	Cin=> '0'	,
	Cout=> Carry( 	2304	),
	S=> R(	37	));
			
  U2305	: Soma_AMA3_1 PORT MAP(
	A=> C(	2369	),
	B=>E(	2206	),
	Cin=> Carry( 	2304	),
	Cout=> Carry( 	2305	),
	S=> E(	2268	));
			
  U2306	: Soma_AMA3_1 PORT MAP(
	A=> C(	2370	),
	B=>E(	2207	),
	Cin=> Carry( 	2305	),
	Cout=> Carry( 	2306	),
	S=> E(	2269	));
			
  U2307	: Soma_AMA3_1 PORT MAP(
	A=> C(	2371	),
	B=>E(	2208	),
	Cin=> Carry( 	2306	),
	Cout=> Carry( 	2307	),
	S=> E(	2270	));
			
  U2308	: Soma_AMA3_1 PORT MAP(
	A=> C(	2372	),
	B=>E(	2209	),
	Cin=> Carry( 	2307	),
	Cout=> Carry( 	2308	),
	S=> E(	2271	));
			
  U2309	: Soma_AMA3_1 PORT MAP(
	A=> C(	2373	),
	B=>E(	2210	),
	Cin=> Carry( 	2308	),
	Cout=> Carry( 	2309	),
	S=> E(	2272	));
			
  U2310	: Soma_AMA3_1 PORT MAP(
	A=> C(	2374	),
	B=>E(	2211	),
	Cin=> Carry( 	2309	),
	Cout=> Carry( 	2310	),
	S=> E(	2273	));
			
  U2311	: Soma_AMA3_1 PORT MAP(
	A=> C(	2375	),
	B=>E(	2212	),
	Cin=> Carry( 	2310	),
	Cout=> Carry( 	2311	),
	S=> E(	2274	));
			
  U2312	: Soma_AMA3_1 PORT MAP(
	A=> C(	2376	),
	B=>E(	2213	),
	Cin=> Carry( 	2311	),
	Cout=> Carry( 	2312	),
	S=> E(	2275	));
			
  U2313	: Soma_AMA3_1 PORT MAP(
	A=> C(	2377	),
	B=>E(	2214	),
	Cin=> Carry( 	2312	),
	Cout=> Carry( 	2313	),
	S=> E(	2276	));
			
  U2314	: Soma_AMA3_1 PORT MAP(
	A=> C(	2378	),
	B=>E(	2215	),
	Cin=> Carry( 	2313	),
	Cout=> Carry( 	2314	),
	S=> E(	2277	));
			
  U2315	: Soma_AMA3_1 PORT MAP(
	A=> C(	2379	),
	B=>E(	2216	),
	Cin=> Carry( 	2314	),
	Cout=> Carry( 	2315	),
	S=> E(	2278	));
			
  U2316	: Soma_AMA3_1 PORT MAP(
	A=> C(	2380	),
	B=>E(	2217	),
	Cin=> Carry( 	2315	),
	Cout=> Carry( 	2316	),
	S=> E(	2279	));
			
  U2317	: Soma_AMA3_1 PORT MAP(
	A=> C(	2381	),
	B=>E(	2218	),
	Cin=> Carry( 	2316	),
	Cout=> Carry( 	2317	),
	S=> E(	2280	));
			
  U2318	: Soma_AMA3_1 PORT MAP(
	A=> C(	2382	),
	B=>E(	2219	),
	Cin=> Carry( 	2317	),
	Cout=> Carry( 	2318	),
	S=> E(	2281	));
			
  U2319	: Soma_AMA3_1 PORT MAP(
	A=> C(	2383	),
	B=>E(	2220	),
	Cin=> Carry( 	2318	),
	Cout=> Carry( 	2319	),
	S=> E(	2282	));
			
  U2320	: Soma_AMA3_1 PORT MAP(
	A=> C(	2384	),
	B=>E(	2221	),
	Cin=> Carry( 	2319	),
	Cout=> Carry( 	2320	),
	S=> E(	2283	));
			
  U2321	: Soma_AMA3_1 PORT MAP(
	A=> C(	2385	),
	B=>E(	2222	),
	Cin=> Carry( 	2320	),
	Cout=> Carry( 	2321	),
	S=> E(	2284	));
			
  U2322	: Soma_AMA3_1 PORT MAP(
	A=> C(	2386	),
	B=>E(	2223	),
	Cin=> Carry( 	2321	),
	Cout=> Carry( 	2322	),
	S=> E(	2285	));
			
  U2323	: Soma_AMA3_1 PORT MAP(
	A=> C(	2387	),
	B=>E(	2224	),
	Cin=> Carry( 	2322	),
	Cout=> Carry( 	2323	),
	S=> E(	2286	));
			
  U2324	: Soma_AMA3_1 PORT MAP(
	A=> C(	2388	),
	B=>E(	2225	),
	Cin=> Carry( 	2323	),
	Cout=> Carry( 	2324	),
	S=> E(	2287	));
			
  U2325	: Soma_AMA3_1 PORT MAP(
	A=> C(	2389	),
	B=>E(	2226	),
	Cin=> Carry( 	2324	),
	Cout=> Carry( 	2325	),
	S=> E(	2288	));
			
  U2326	: Soma_AMA3_1 PORT MAP(
	A=> C(	2390	),
	B=>E(	2227	),
	Cin=> Carry( 	2325	),
	Cout=> Carry( 	2326	),
	S=> E(	2289	));
			
  U2327	: Soma_AMA3_1 PORT MAP(
	A=> C(	2391	),
	B=>E(	2228	),
	Cin=> Carry( 	2326	),
	Cout=> Carry( 	2327	),
	S=> E(	2290	));
			
  U2328	: Soma_AMA3_1 PORT MAP(
	A=> C(	2392	),
	B=>E(	2229	),
	Cin=> Carry( 	2327	),
	Cout=> Carry( 	2328	),
	S=> E(	2291	));
			
  U2329	: Soma_AMA3_1 PORT MAP(
	A=> C(	2393	),
	B=>E(	2230	),
	Cin=> Carry( 	2328	),
	Cout=> Carry( 	2329	),
	S=> E(	2292	));
			
  U2330	: Soma_AMA3_1 PORT MAP(
	A=> C(	2394	),
	B=>E(	2231	),
	Cin=> Carry( 	2329	),
	Cout=> Carry( 	2330	),
	S=> E(	2293	));
			
  U2331	: Soma_AMA3_1 PORT MAP(
	A=> C(	2395	),
	B=>E(	2232	),
	Cin=> Carry( 	2330	),
	Cout=> Carry( 	2331	),
	S=> E(	2294	));
			
  U2332	: Soma_AMA3_1 PORT MAP(
	A=> C(	2396	),
	B=>E(	2233	),
	Cin=> Carry( 	2331	),
	Cout=> Carry( 	2332	),
	S=> E(	2295	));
			
  U2333	: Soma_AMA3_1 PORT MAP(
	A=> C(	2397	),
	B=>E(	2234	),
	Cin=> Carry( 	2332	),
	Cout=> Carry( 	2333	),
	S=> E(	2296	));
			
  U2334	: Soma_AMA3_1 PORT MAP(
	A=> C(	2398	),
	B=>E(	2235	),
	Cin=> Carry( 	2333	),
	Cout=> Carry( 	2334	),
	S=> E(	2297	));
			
  U2335	: Soma_AMA3_1 PORT MAP(
	A=> C(	2399	),
	B=>E(	2236	),
	Cin=> Carry( 	2334	),
	Cout=> Carry( 	2335	),
	S=> E(	2298	));
			
  U2336	: Soma_AMA3_1 PORT MAP(
	A=> C(	2400	),
	B=>E(	2237	),
	Cin=> Carry( 	2335	),
	Cout=> Carry( 	2336	),
	S=> E(	2299	));
			
  U2337	: Soma_AMA3_1 PORT MAP(
	A=> C(	2401	),
	B=>E(	2238	),
	Cin=> Carry( 	2336	),
	Cout=> Carry( 	2337	),
	S=> E(	2300	));
			
  U2338	: Soma_AMA3_1 PORT MAP(
	A=> C(	2402	),
	B=>E(	2239	),
	Cin=> Carry( 	2337	),
	Cout=> Carry( 	2338	),
	S=> E(	2301	));
			
  U2339	: Soma_AMA3_1 PORT MAP(
	A=> C(	2403	),
	B=>E(	2240	),
	Cin=> Carry( 	2338	),
	Cout=> Carry( 	2339	),
	S=> E(	2302	));
			
  U2340	: Soma_AMA3_1 PORT MAP(
	A=> C(	2404	),
	B=>E(	2241	),
	Cin=> Carry( 	2339	),
	Cout=> Carry( 	2340	),
	S=> E(	2303	));
			
  U2341	: Soma_AMA3_1 PORT MAP(
	A=> C(	2405	),
	B=>E(	2242	),
	Cin=> Carry( 	2340	),
	Cout=> Carry( 	2341	),
	S=> E(	2304	));
			
  U2342	: Soma_AMA3_1 PORT MAP(
	A=> C(	2406	),
	B=>E(	2243	),
	Cin=> Carry( 	2341	),
	Cout=> Carry( 	2342	),
	S=> E(	2305	));
			
  U2343	: Soma_AMA3_1 PORT MAP(
	A=> C(	2407	),
	B=>E(	2244	),
	Cin=> Carry( 	2342	),
	Cout=> Carry( 	2343	),
	S=> E(	2306	));
			
  U2344	: Soma_AMA3_1 PORT MAP(
	A=> C(	2408	),
	B=>E(	2245	),
	Cin=> Carry( 	2343	),
	Cout=> Carry( 	2344	),
	S=> E(	2307	));
			
  U2345	: Soma_AMA3_1 PORT MAP(
	A=> C(	2409	),
	B=>E(	2246	),
	Cin=> Carry( 	2344	),
	Cout=> Carry( 	2345	),
	S=> E(	2308	));
			
  U2346	: Soma_AMA3_1 PORT MAP(
	A=> C(	2410	),
	B=>E(	2247	),
	Cin=> Carry( 	2345	),
	Cout=> Carry( 	2346	),
	S=> E(	2309	));
			
  U2347	: Soma_AMA3_1 PORT MAP(
	A=> C(	2411	),
	B=>E(	2248	),
	Cin=> Carry( 	2346	),
	Cout=> Carry( 	2347	),
	S=> E(	2310	));
			
  U2348	: Soma_AMA3_1 PORT MAP(
	A=> C(	2412	),
	B=>E(	2249	),
	Cin=> Carry( 	2347	),
	Cout=> Carry( 	2348	),
	S=> E(	2311	));
			
  U2349	: Soma_AMA3_1 PORT MAP(
	A=> C(	2413	),
	B=>E(	2250	),
	Cin=> Carry( 	2348	),
	Cout=> Carry( 	2349	),
	S=> E(	2312	));
			
  U2350	: Soma_AMA3_1 PORT MAP(
	A=> C(	2414	),
	B=>E(	2251	),
	Cin=> Carry( 	2349	),
	Cout=> Carry( 	2350	),
	S=> E(	2313	));
			
  U2351	: Soma_AMA3_1 PORT MAP(
	A=> C(	2415	),
	B=>E(	2252	),
	Cin=> Carry( 	2350	),
	Cout=> Carry( 	2351	),
	S=> E(	2314	));
			
  U2352	: Soma_AMA3_1 PORT MAP(
	A=> C(	2416	),
	B=>E(	2253	),
	Cin=> Carry( 	2351	),
	Cout=> Carry( 	2352	),
	S=> E(	2315	));
			
  U2353	: Soma_AMA3_1 PORT MAP(
	A=> C(	2417	),
	B=>E(	2254	),
	Cin=> Carry( 	2352	),
	Cout=> Carry( 	2353	),
	S=> E(	2316	));
			
  U2354	: Soma_AMA3_1 PORT MAP(
	A=> C(	2418	),
	B=>E(	2255	),
	Cin=> Carry( 	2353	),
	Cout=> Carry( 	2354	),
	S=> E(	2317	));
			
  U2355	: Soma_AMA3_1 PORT MAP(
	A=> C(	2419	),
	B=>E(	2256	),
	Cin=> Carry( 	2354	),
	Cout=> Carry( 	2355	),
	S=> E(	2318	));
			
  U2356	: Soma_AMA3_1 PORT MAP(
	A=> C(	2420	),
	B=>E(	2257	),
	Cin=> Carry( 	2355	),
	Cout=> Carry( 	2356	),
	S=> E(	2319	));
			
  U2357	: Soma_AMA3_1 PORT MAP(
	A=> C(	2421	),
	B=>E(	2258	),
	Cin=> Carry( 	2356	),
	Cout=> Carry( 	2357	),
	S=> E(	2320	));
			
  U2358	: Soma_AMA3_1 PORT MAP(
	A=> C(	2422	),
	B=>E(	2259	),
	Cin=> Carry( 	2357	),
	Cout=> Carry( 	2358	),
	S=> E(	2321	));
			
  U2359	: Soma_AMA3_1 PORT MAP(
	A=> C(	2423	),
	B=>E(	2260	),
	Cin=> Carry( 	2358	),
	Cout=> Carry( 	2359	),
	S=> E(	2322	));
			
  U2360	: Soma_AMA3_1 PORT MAP(
	A=> C(	2424	),
	B=>E(	2261	),
	Cin=> Carry( 	2359	),
	Cout=> Carry( 	2360	),
	S=> E(	2323	));
			
  U2361	: Soma_AMA3_1 PORT MAP(
	A=> C(	2425	),
	B=>E(	2262	),
	Cin=> Carry( 	2360	),
	Cout=> Carry( 	2361	),
	S=> E(	2324	));
			
  U2362	: Soma_AMA3_1 PORT MAP(
	A=> C(	2426	),
	B=>E(	2263	),
	Cin=> Carry( 	2361	),
	Cout=> Carry( 	2362	),
	S=> E(	2325	));
			
  U2363	: Soma_AMA3_1 PORT MAP(
	A=> C(	2427	),
	B=>E(	2264	),
	Cin=> Carry( 	2362	),
	Cout=> Carry( 	2363	),
	S=> E(	2326	));
			
  U2364	: Soma_AMA3_1 PORT MAP(
	A=> C(	2428	),
	B=>E(	2265	),
	Cin=> Carry( 	2363	),
	Cout=> Carry( 	2364	),
	S=> E(	2327	));
			
  U2365	: Soma_AMA3_1 PORT MAP(
	A=> C(	2429	),
	B=>E(	2266	),
	Cin=> Carry( 	2364	),
	Cout=> Carry( 	2365	),
	S=> E(	2328	));
			
  U2366	: Soma_AMA3_1 PORT MAP(
	A=> C(	2430	),
	B=>E(	2267	),
	Cin=> Carry( 	2365	),
	Cout=> Carry( 	2366	),
	S=> E(	2329	));
			
U2367	: Soma_AMA3_1 PORT MAP(
	A=> C(	2431	),
	B=>Carry(	2303	),
	Cin=> Carry( 	2366	),
	Cout=> Carry( 	2367	),
	S=> E(	2330	));

			
  U2368	: Soma_AMA3_1 PORT MAP(
	A=> C(	2432	),
	B=>E(	2268	),
	Cin=> '0'	,
	Cout=> Carry( 	2368	),
	S=> R(	38	));
			
  U2369	: Soma_AMA3_1 PORT MAP(
	A=> C(	2433	),
	B=>E(	2269	),
	Cin=> Carry( 	2368	),
	Cout=> Carry( 	2369	),
	S=> E(	2331	));
			
  U2370	: Soma_AMA3_1 PORT MAP(
	A=> C(	2434	),
	B=>E(	2270	),
	Cin=> Carry( 	2369	),
	Cout=> Carry( 	2370	),
	S=> E(	2332	));
			
  U2371	: Soma_AMA3_1 PORT MAP(
	A=> C(	2435	),
	B=>E(	2271	),
	Cin=> Carry( 	2370	),
	Cout=> Carry( 	2371	),
	S=> E(	2333	));
			
  U2372	: Soma_AMA3_1 PORT MAP(
	A=> C(	2436	),
	B=>E(	2272	),
	Cin=> Carry( 	2371	),
	Cout=> Carry( 	2372	),
	S=> E(	2334	));
			
  U2373	: Soma_AMA3_1 PORT MAP(
	A=> C(	2437	),
	B=>E(	2273	),
	Cin=> Carry( 	2372	),
	Cout=> Carry( 	2373	),
	S=> E(	2335	));
			
  U2374	: Soma_AMA3_1 PORT MAP(
	A=> C(	2438	),
	B=>E(	2274	),
	Cin=> Carry( 	2373	),
	Cout=> Carry( 	2374	),
	S=> E(	2336	));
			
  U2375	: Soma_AMA3_1 PORT MAP(
	A=> C(	2439	),
	B=>E(	2275	),
	Cin=> Carry( 	2374	),
	Cout=> Carry( 	2375	),
	S=> E(	2337	));
			
  U2376	: Soma_AMA3_1 PORT MAP(
	A=> C(	2440	),
	B=>E(	2276	),
	Cin=> Carry( 	2375	),
	Cout=> Carry( 	2376	),
	S=> E(	2338	));
			
  U2377	: Soma_AMA3_1 PORT MAP(
	A=> C(	2441	),
	B=>E(	2277	),
	Cin=> Carry( 	2376	),
	Cout=> Carry( 	2377	),
	S=> E(	2339	));
			
  U2378	: Soma_AMA3_1 PORT MAP(
	A=> C(	2442	),
	B=>E(	2278	),
	Cin=> Carry( 	2377	),
	Cout=> Carry( 	2378	),
	S=> E(	2340	));
			
  U2379	: Soma_AMA3_1 PORT MAP(
	A=> C(	2443	),
	B=>E(	2279	),
	Cin=> Carry( 	2378	),
	Cout=> Carry( 	2379	),
	S=> E(	2341	));
			
  U2380	: Soma_AMA3_1 PORT MAP(
	A=> C(	2444	),
	B=>E(	2280	),
	Cin=> Carry( 	2379	),
	Cout=> Carry( 	2380	),
	S=> E(	2342	));
			
  U2381	: Soma_AMA3_1 PORT MAP(
	A=> C(	2445	),
	B=>E(	2281	),
	Cin=> Carry( 	2380	),
	Cout=> Carry( 	2381	),
	S=> E(	2343	));
			
  U2382	: Soma_AMA3_1 PORT MAP(
	A=> C(	2446	),
	B=>E(	2282	),
	Cin=> Carry( 	2381	),
	Cout=> Carry( 	2382	),
	S=> E(	2344	));
			
  U2383	: Soma_AMA3_1 PORT MAP(
	A=> C(	2447	),
	B=>E(	2283	),
	Cin=> Carry( 	2382	),
	Cout=> Carry( 	2383	),
	S=> E(	2345	));
			
  U2384	: Soma_AMA3_1 PORT MAP(
	A=> C(	2448	),
	B=>E(	2284	),
	Cin=> Carry( 	2383	),
	Cout=> Carry( 	2384	),
	S=> E(	2346	));
			
  U2385	: Soma_AMA3_1 PORT MAP(
	A=> C(	2449	),
	B=>E(	2285	),
	Cin=> Carry( 	2384	),
	Cout=> Carry( 	2385	),
	S=> E(	2347	));
			
  U2386	: Soma_AMA3_1 PORT MAP(
	A=> C(	2450	),
	B=>E(	2286	),
	Cin=> Carry( 	2385	),
	Cout=> Carry( 	2386	),
	S=> E(	2348	));
			
  U2387	: Soma_AMA3_1 PORT MAP(
	A=> C(	2451	),
	B=>E(	2287	),
	Cin=> Carry( 	2386	),
	Cout=> Carry( 	2387	),
	S=> E(	2349	));
			
  U2388	: Soma_AMA3_1 PORT MAP(
	A=> C(	2452	),
	B=>E(	2288	),
	Cin=> Carry( 	2387	),
	Cout=> Carry( 	2388	),
	S=> E(	2350	));
			
  U2389	: Soma_AMA3_1 PORT MAP(
	A=> C(	2453	),
	B=>E(	2289	),
	Cin=> Carry( 	2388	),
	Cout=> Carry( 	2389	),
	S=> E(	2351	));
			
  U2390	: Soma_AMA3_1 PORT MAP(
	A=> C(	2454	),
	B=>E(	2290	),
	Cin=> Carry( 	2389	),
	Cout=> Carry( 	2390	),
	S=> E(	2352	));
			
  U2391	: Soma_AMA3_1 PORT MAP(
	A=> C(	2455	),
	B=>E(	2291	),
	Cin=> Carry( 	2390	),
	Cout=> Carry( 	2391	),
	S=> E(	2353	));
			
  U2392	: Soma_AMA3_1 PORT MAP(
	A=> C(	2456	),
	B=>E(	2292	),
	Cin=> Carry( 	2391	),
	Cout=> Carry( 	2392	),
	S=> E(	2354	));
			
  U2393	: Soma_AMA3_1 PORT MAP(
	A=> C(	2457	),
	B=>E(	2293	),
	Cin=> Carry( 	2392	),
	Cout=> Carry( 	2393	),
	S=> E(	2355	));
			
  U2394	: Soma_AMA3_1 PORT MAP(
	A=> C(	2458	),
	B=>E(	2294	),
	Cin=> Carry( 	2393	),
	Cout=> Carry( 	2394	),
	S=> E(	2356	));
			
  U2395	: Soma_AMA3_1 PORT MAP(
	A=> C(	2459	),
	B=>E(	2295	),
	Cin=> Carry( 	2394	),
	Cout=> Carry( 	2395	),
	S=> E(	2357	));
			
  U2396	: Soma_AMA3_1 PORT MAP(
	A=> C(	2460	),
	B=>E(	2296	),
	Cin=> Carry( 	2395	),
	Cout=> Carry( 	2396	),
	S=> E(	2358	));
			
  U2397	: Soma_AMA3_1 PORT MAP(
	A=> C(	2461	),
	B=>E(	2297	),
	Cin=> Carry( 	2396	),
	Cout=> Carry( 	2397	),
	S=> E(	2359	));
			
  U2398	: Soma_AMA3_1 PORT MAP(
	A=> C(	2462	),
	B=>E(	2298	),
	Cin=> Carry( 	2397	),
	Cout=> Carry( 	2398	),
	S=> E(	2360	));
			
  U2399	: Soma_AMA3_1 PORT MAP(
	A=> C(	2463	),
	B=>E(	2299	),
	Cin=> Carry( 	2398	),
	Cout=> Carry( 	2399	),
	S=> E(	2361	));
			
  U2400	: Soma_AMA3_1 PORT MAP(
	A=> C(	2464	),
	B=>E(	2300	),
	Cin=> Carry( 	2399	),
	Cout=> Carry( 	2400	),
	S=> E(	2362	));
			
  U2401	: Soma_AMA3_1 PORT MAP(
	A=> C(	2465	),
	B=>E(	2301	),
	Cin=> Carry( 	2400	),
	Cout=> Carry( 	2401	),
	S=> E(	2363	));
			
  U2402	: Soma_AMA3_1 PORT MAP(
	A=> C(	2466	),
	B=>E(	2302	),
	Cin=> Carry( 	2401	),
	Cout=> Carry( 	2402	),
	S=> E(	2364	));
			
  U2403	: Soma_AMA3_1 PORT MAP(
	A=> C(	2467	),
	B=>E(	2303	),
	Cin=> Carry( 	2402	),
	Cout=> Carry( 	2403	),
	S=> E(	2365	));
			
  U2404	: Soma_AMA3_1 PORT MAP(
	A=> C(	2468	),
	B=>E(	2304	),
	Cin=> Carry( 	2403	),
	Cout=> Carry( 	2404	),
	S=> E(	2366	));
			
  U2405	: Soma_AMA3_1 PORT MAP(
	A=> C(	2469	),
	B=>E(	2305	),
	Cin=> Carry( 	2404	),
	Cout=> Carry( 	2405	),
	S=> E(	2367	));
			
  U2406	: Soma_AMA3_1 PORT MAP(
	A=> C(	2470	),
	B=>E(	2306	),
	Cin=> Carry( 	2405	),
	Cout=> Carry( 	2406	),
	S=> E(	2368	));
			
  U2407	: Soma_AMA3_1 PORT MAP(
	A=> C(	2471	),
	B=>E(	2307	),
	Cin=> Carry( 	2406	),
	Cout=> Carry( 	2407	),
	S=> E(	2369	));
			
  U2408	: Soma_AMA3_1 PORT MAP(
	A=> C(	2472	),
	B=>E(	2308	),
	Cin=> Carry( 	2407	),
	Cout=> Carry( 	2408	),
	S=> E(	2370	));
			
  U2409	: Soma_AMA3_1 PORT MAP(
	A=> C(	2473	),
	B=>E(	2309	),
	Cin=> Carry( 	2408	),
	Cout=> Carry( 	2409	),
	S=> E(	2371	));
			
  U2410	: Soma_AMA3_1 PORT MAP(
	A=> C(	2474	),
	B=>E(	2310	),
	Cin=> Carry( 	2409	),
	Cout=> Carry( 	2410	),
	S=> E(	2372	));
			
  U2411	: Soma_AMA3_1 PORT MAP(
	A=> C(	2475	),
	B=>E(	2311	),
	Cin=> Carry( 	2410	),
	Cout=> Carry( 	2411	),
	S=> E(	2373	));
			
  U2412	: Soma_AMA3_1 PORT MAP(
	A=> C(	2476	),
	B=>E(	2312	),
	Cin=> Carry( 	2411	),
	Cout=> Carry( 	2412	),
	S=> E(	2374	));
			
  U2413	: Soma_AMA3_1 PORT MAP(
	A=> C(	2477	),
	B=>E(	2313	),
	Cin=> Carry( 	2412	),
	Cout=> Carry( 	2413	),
	S=> E(	2375	));
			
  U2414	: Soma_AMA3_1 PORT MAP(
	A=> C(	2478	),
	B=>E(	2314	),
	Cin=> Carry( 	2413	),
	Cout=> Carry( 	2414	),
	S=> E(	2376	));
			
  U2415	: Soma_AMA3_1 PORT MAP(
	A=> C(	2479	),
	B=>E(	2315	),
	Cin=> Carry( 	2414	),
	Cout=> Carry( 	2415	),
	S=> E(	2377	));
			
  U2416	: Soma_AMA3_1 PORT MAP(
	A=> C(	2480	),
	B=>E(	2316	),
	Cin=> Carry( 	2415	),
	Cout=> Carry( 	2416	),
	S=> E(	2378	));
			
  U2417	: Soma_AMA3_1 PORT MAP(
	A=> C(	2481	),
	B=>E(	2317	),
	Cin=> Carry( 	2416	),
	Cout=> Carry( 	2417	),
	S=> E(	2379	));
			
  U2418	: Soma_AMA3_1 PORT MAP(
	A=> C(	2482	),
	B=>E(	2318	),
	Cin=> Carry( 	2417	),
	Cout=> Carry( 	2418	),
	S=> E(	2380	));
			
  U2419	: Soma_AMA3_1 PORT MAP(
	A=> C(	2483	),
	B=>E(	2319	),
	Cin=> Carry( 	2418	),
	Cout=> Carry( 	2419	),
	S=> E(	2381	));
			
  U2420	: Soma_AMA3_1 PORT MAP(
	A=> C(	2484	),
	B=>E(	2320	),
	Cin=> Carry( 	2419	),
	Cout=> Carry( 	2420	),
	S=> E(	2382	));
			
  U2421	: Soma_AMA3_1 PORT MAP(
	A=> C(	2485	),
	B=>E(	2321	),
	Cin=> Carry( 	2420	),
	Cout=> Carry( 	2421	),
	S=> E(	2383	));
			
  U2422	: Soma_AMA3_1 PORT MAP(
	A=> C(	2486	),
	B=>E(	2322	),
	Cin=> Carry( 	2421	),
	Cout=> Carry( 	2422	),
	S=> E(	2384	));
			
  U2423	: Soma_AMA3_1 PORT MAP(
	A=> C(	2487	),
	B=>E(	2323	),
	Cin=> Carry( 	2422	),
	Cout=> Carry( 	2423	),
	S=> E(	2385	));
			
  U2424	: Soma_AMA3_1 PORT MAP(
	A=> C(	2488	),
	B=>E(	2324	),
	Cin=> Carry( 	2423	),
	Cout=> Carry( 	2424	),
	S=> E(	2386	));
			
  U2425	: Soma_AMA3_1 PORT MAP(
	A=> C(	2489	),
	B=>E(	2325	),
	Cin=> Carry( 	2424	),
	Cout=> Carry( 	2425	),
	S=> E(	2387	));
			
  U2426	: Soma_AMA3_1 PORT MAP(
	A=> C(	2490	),
	B=>E(	2326	),
	Cin=> Carry( 	2425	),
	Cout=> Carry( 	2426	),
	S=> E(	2388	));
			
  U2427	: Soma_AMA3_1 PORT MAP(
	A=> C(	2491	),
	B=>E(	2327	),
	Cin=> Carry( 	2426	),
	Cout=> Carry( 	2427	),
	S=> E(	2389	));
			
  U2428	: Soma_AMA3_1 PORT MAP(
	A=> C(	2492	),
	B=>E(	2328	),
	Cin=> Carry( 	2427	),
	Cout=> Carry( 	2428	),
	S=> E(	2390	));
			
  U2429	: Soma_AMA3_1 PORT MAP(
	A=> C(	2493	),
	B=>E(	2329	),
	Cin=> Carry( 	2428	),
	Cout=> Carry( 	2429	),
	S=> E(	2391	));
			
  U2430	: Soma_AMA3_1 PORT MAP(
	A=> C(	2494	),
	B=>E(	2330	),
	Cin=> Carry( 	2429	),
	Cout=> Carry( 	2430	),
	S=> E(	2392	));
			
  U2431	: Soma_AMA3_1 PORT MAP(
	A=> C(	2495	),
	B=>Carry(	2367	),
	Cin=> Carry( 	2430	),
	Cout=> Carry( 	2431	),
	S=> E(	2393	));

			
  U2432	: Soma_AMA3_1 PORT MAP(
	A=> C(	2496	),
	B=>E(	2331	),
	Cin=>'0'	,
	Cout=> Carry( 	2432	),
	S=> R(	39	));
			
  U2433	: Soma_AMA3_1 PORT MAP(
	A=> C(	2497	),
	B=>E(	2332	),
	Cin=> Carry( 	2432	),
	Cout=> Carry( 	2433	),
	S=> E(	2394	));
			
  U2434	: Soma_AMA3_1 PORT MAP(
	A=> C(	2498	),
	B=>E(	2333	),
	Cin=> Carry( 	2433	),
	Cout=> Carry( 	2434	),
	S=> E(	2395	));
			
  U2435	: Soma_AMA3_1 PORT MAP(
	A=> C(	2499	),
	B=>E(	2334	),
	Cin=> Carry( 	2434	),
	Cout=> Carry( 	2435	),
	S=> E(	2396	));
			
  U2436	: Soma_AMA3_1 PORT MAP(
	A=> C(	2500	),
	B=>E(	2335	),
	Cin=> Carry( 	2435	),
	Cout=> Carry( 	2436	),
	S=> E(	2397	));
			
  U2437	: Soma_AMA3_1 PORT MAP(
	A=> C(	2501	),
	B=>E(	2336	),
	Cin=> Carry( 	2436	),
	Cout=> Carry( 	2437	),
	S=> E(	2398	));
			
  U2438	: Soma_AMA3_1 PORT MAP(
	A=> C(	2502	),
	B=>E(	2337	),
	Cin=> Carry( 	2437	),
	Cout=> Carry( 	2438	),
	S=> E(	2399	));
			
  U2439	: Soma_AMA3_1 PORT MAP(
	A=> C(	2503	),
	B=>E(	2338	),
	Cin=> Carry( 	2438	),
	Cout=> Carry( 	2439	),
	S=> E(	2400	));
			
  U2440	: Soma_AMA3_1 PORT MAP(
	A=> C(	2504	),
	B=>E(	2339	),
	Cin=> Carry( 	2439	),
	Cout=> Carry( 	2440	),
	S=> E(	2401	));
			
  U2441	: Soma_AMA3_1 PORT MAP(
	A=> C(	2505	),
	B=>E(	2340	),
	Cin=> Carry( 	2440	),
	Cout=> Carry( 	2441	),
	S=> E(	2402	));
			
  U2442	: Soma_AMA3_1 PORT MAP(
	A=> C(	2506	),
	B=>E(	2341	),
	Cin=> Carry( 	2441	),
	Cout=> Carry( 	2442	),
	S=> E(	2403	));
			
  U2443	: Soma_AMA3_1 PORT MAP(
	A=> C(	2507	),
	B=>E(	2342	),
	Cin=> Carry( 	2442	),
	Cout=> Carry( 	2443	),
	S=> E(	2404	));
			
  U2444	: Soma_AMA3_1 PORT MAP(
	A=> C(	2508	),
	B=>E(	2343	),
	Cin=> Carry( 	2443	),
	Cout=> Carry( 	2444	),
	S=> E(	2405	));
			
  U2445	: Soma_AMA3_1 PORT MAP(
	A=> C(	2509	),
	B=>E(	2344	),
	Cin=> Carry( 	2444	),
	Cout=> Carry( 	2445	),
	S=> E(	2406	));
			
  U2446	: Soma_AMA3_1 PORT MAP(
	A=> C(	2510	),
	B=>E(	2345	),
	Cin=> Carry( 	2445	),
	Cout=> Carry( 	2446	),
	S=> E(	2407	));
			
  U2447	: Soma_AMA3_1 PORT MAP(
	A=> C(	2511	),
	B=>E(	2346	),
	Cin=> Carry( 	2446	),
	Cout=> Carry( 	2447	),
	S=> E(	2408	));
			
  U2448	: Soma_AMA3_1 PORT MAP(
	A=> C(	2512	),
	B=>E(	2347	),
	Cin=> Carry( 	2447	),
	Cout=> Carry( 	2448	),
	S=> E(	2409	));
			
  U2449	: Soma_AMA3_1 PORT MAP(
	A=> C(	2513	),
	B=>E(	2348	),
	Cin=> Carry( 	2448	),
	Cout=> Carry( 	2449	),
	S=> E(	2410	));
			
  U2450	: Soma_AMA3_1 PORT MAP(
	A=> C(	2514	),
	B=>E(	2349	),
	Cin=> Carry( 	2449	),
	Cout=> Carry( 	2450	),
	S=> E(	2411	));
			
  U2451	: Soma_AMA3_1 PORT MAP(
	A=> C(	2515	),
	B=>E(	2350	),
	Cin=> Carry( 	2450	),
	Cout=> Carry( 	2451	),
	S=> E(	2412	));
			
  U2452	: Soma_AMA3_1 PORT MAP(
	A=> C(	2516	),
	B=>E(	2351	),
	Cin=> Carry( 	2451	),
	Cout=> Carry( 	2452	),
	S=> E(	2413	));
			
  U2453	: Soma_AMA3_1 PORT MAP(
	A=> C(	2517	),
	B=>E(	2352	),
	Cin=> Carry( 	2452	),
	Cout=> Carry( 	2453	),
	S=> E(	2414	));
			
  U2454	: Soma_AMA3_1 PORT MAP(
	A=> C(	2518	),
	B=>E(	2353	),
	Cin=> Carry( 	2453	),
	Cout=> Carry( 	2454	),
	S=> E(	2415	));
			
  U2455	: Soma_AMA3_1 PORT MAP(
	A=> C(	2519	),
	B=>E(	2354	),
	Cin=> Carry( 	2454	),
	Cout=> Carry( 	2455	),
	S=> E(	2416	));
			
  U2456	: Soma_AMA3_1 PORT MAP(
	A=> C(	2520	),
	B=>E(	2355	),
	Cin=> Carry( 	2455	),
	Cout=> Carry( 	2456	),
	S=> E(	2417	));
			
  U2457	: Soma_AMA3_1 PORT MAP(
	A=> C(	2521	),
	B=>E(	2356	),
	Cin=> Carry( 	2456	),
	Cout=> Carry( 	2457	),
	S=> E(	2418	));
			
  U2458	: Soma_AMA3_1 PORT MAP(
	A=> C(	2522	),
	B=>E(	2357	),
	Cin=> Carry( 	2457	),
	Cout=> Carry( 	2458	),
	S=> E(	2419	));
			
  U2459	: Soma_AMA3_1 PORT MAP(
	A=> C(	2523	),
	B=>E(	2358	),
	Cin=> Carry( 	2458	),
	Cout=> Carry( 	2459	),
	S=> E(	2420	));
			
  U2460	: Soma_AMA3_1 PORT MAP(
	A=> C(	2524	),
	B=>E(	2359	),
	Cin=> Carry( 	2459	),
	Cout=> Carry( 	2460	),
	S=> E(	2421	));
			
  U2461	: Soma_AMA3_1 PORT MAP(
	A=> C(	2525	),
	B=>E(	2360	),
	Cin=> Carry( 	2460	),
	Cout=> Carry( 	2461	),
	S=> E(	2422	));
			
  U2462	: Soma_AMA3_1 PORT MAP(
	A=> C(	2526	),
	B=>E(	2361	),
	Cin=> Carry( 	2461	),
	Cout=> Carry( 	2462	),
	S=> E(	2423	));
			
  U2463	: Soma_AMA3_1 PORT MAP(
	A=> C(	2527	),
	B=>E(	2362	),
	Cin=> Carry( 	2462	),
	Cout=> Carry( 	2463	),
	S=> E(	2424	));
			
  U2464	: Soma_AMA3_1 PORT MAP(
	A=> C(	2528	),
	B=>E(	2363	),
	Cin=> Carry( 	2463	),
	Cout=> Carry( 	2464	),
	S=> E(	2425	));
			
  U2465	: Soma_AMA3_1 PORT MAP(
	A=> C(	2529	),
	B=>E(	2364	),
	Cin=> Carry( 	2464	),
	Cout=> Carry( 	2465	),
	S=> E(	2426	));
			
  U2466	: Soma_AMA3_1 PORT MAP(
	A=> C(	2530	),
	B=>E(	2365	),
	Cin=> Carry( 	2465	),
	Cout=> Carry( 	2466	),
	S=> E(	2427	));
			
  U2467	: Soma_AMA3_1 PORT MAP(
	A=> C(	2531	),
	B=>E(	2366	),
	Cin=> Carry( 	2466	),
	Cout=> Carry( 	2467	),
	S=> E(	2428	));
			
  U2468	: Soma_AMA3_1 PORT MAP(
	A=> C(	2532	),
	B=>E(	2367	),
	Cin=> Carry( 	2467	),
	Cout=> Carry( 	2468	),
	S=> E(	2429	));
			
  U2469	: Soma_AMA3_1 PORT MAP(
	A=> C(	2533	),
	B=>E(	2368	),
	Cin=> Carry( 	2468	),
	Cout=> Carry( 	2469	),
	S=> E(	2430	));
			
  U2470	: Soma_AMA3_1 PORT MAP(
	A=> C(	2534	),
	B=>E(	2369	),
	Cin=> Carry( 	2469	),
	Cout=> Carry( 	2470	),
	S=> E(	2431	));
			
  U2471	: Soma_AMA3_1 PORT MAP(
	A=> C(	2535	),
	B=>E(	2370	),
	Cin=> Carry( 	2470	),
	Cout=> Carry( 	2471	),
	S=> E(	2432	));
			
  U2472	: Soma_AMA3_1 PORT MAP(
	A=> C(	2536	),
	B=>E(	2371	),
	Cin=> Carry( 	2471	),
	Cout=> Carry( 	2472	),
	S=> E(	2433	));
			
  U2473	: Soma_AMA3_1 PORT MAP(
	A=> C(	2537	),
	B=>E(	2372	),
	Cin=> Carry( 	2472	),
	Cout=> Carry( 	2473	),
	S=> E(	2434	));
			
  U2474	: Soma_AMA3_1 PORT MAP(
	A=> C(	2538	),
	B=>E(	2373	),
	Cin=> Carry( 	2473	),
	Cout=> Carry( 	2474	),
	S=> E(	2435	));
			
  U2475	: Soma_AMA3_1 PORT MAP(
	A=> C(	2539	),
	B=>E(	2374	),
	Cin=> Carry( 	2474	),
	Cout=> Carry( 	2475	),
	S=> E(	2436	));
			
  U2476	: Soma_AMA3_1 PORT MAP(
	A=> C(	2540	),
	B=>E(	2375	),
	Cin=> Carry( 	2475	),
	Cout=> Carry( 	2476	),
	S=> E(	2437	));
			
  U2477	: Soma_AMA3_1 PORT MAP(
	A=> C(	2541	),
	B=>E(	2376	),
	Cin=> Carry( 	2476	),
	Cout=> Carry( 	2477	),
	S=> E(	2438	));
			
  U2478	: Soma_AMA3_1 PORT MAP(
	A=> C(	2542	),
	B=>E(	2377	),
	Cin=> Carry( 	2477	),
	Cout=> Carry( 	2478	),
	S=> E(	2439	));
			
  U2479	: Soma_AMA3_1 PORT MAP(
	A=> C(	2543	),
	B=>E(	2378	),
	Cin=> Carry( 	2478	),
	Cout=> Carry( 	2479	),
	S=> E(	2440	));
			
  U2480	: Soma_AMA3_1 PORT MAP(
	A=> C(	2544	),
	B=>E(	2379	),
	Cin=> Carry( 	2479	),
	Cout=> Carry( 	2480	),
	S=> E(	2441	));
			
  U2481	: Soma_AMA3_1 PORT MAP(
	A=> C(	2545	),
	B=>E(	2380	),
	Cin=> Carry( 	2480	),
	Cout=> Carry( 	2481	),
	S=> E(	2442	));
			
  U2482	: Soma_AMA3_1 PORT MAP(
	A=> C(	2546	),
	B=>E(	2381	),
	Cin=> Carry( 	2481	),
	Cout=> Carry( 	2482	),
	S=> E(	2443	));
			
  U2483	: Soma_AMA3_1 PORT MAP(
	A=> C(	2547	),
	B=>E(	2382	),
	Cin=> Carry( 	2482	),
	Cout=> Carry( 	2483	),
	S=> E(	2444	));
			
  U2484	: Soma_AMA3_1 PORT MAP(
	A=> C(	2548	),
	B=>E(	2383	),
	Cin=> Carry( 	2483	),
	Cout=> Carry( 	2484	),
	S=> E(	2445	));
			
  U2485	: Soma_AMA3_1 PORT MAP(
	A=> C(	2549	),
	B=>E(	2384	),
	Cin=> Carry( 	2484	),
	Cout=> Carry( 	2485	),
	S=> E(	2446	));
			
  U2486	: Soma_AMA3_1 PORT MAP(
	A=> C(	2550	),
	B=>E(	2385	),
	Cin=> Carry( 	2485	),
	Cout=> Carry( 	2486	),
	S=> E(	2447	));
			
  U2487	: Soma_AMA3_1 PORT MAP(
	A=> C(	2551	),
	B=>E(	2386	),
	Cin=> Carry( 	2486	),
	Cout=> Carry( 	2487	),
	S=> E(	2448	));
			
  U2488	: Soma_AMA3_1 PORT MAP(
	A=> C(	2552	),
	B=>E(	2387	),
	Cin=> Carry( 	2487	),
	Cout=> Carry( 	2488	),
	S=> E(	2449	));
			
  U2489	: Soma_AMA3_1 PORT MAP(
	A=> C(	2553	),
	B=>E(	2388	),
	Cin=> Carry( 	2488	),
	Cout=> Carry( 	2489	),
	S=> E(	2450	));
			
  U2490	: Soma_AMA3_1 PORT MAP(
	A=> C(	2554	),
	B=>E(	2389	),
	Cin=> Carry( 	2489	),
	Cout=> Carry( 	2490	),
	S=> E(	2451	));
			
  U2491	: Soma_AMA3_1 PORT MAP(
	A=> C(	2555	),
	B=>E(	2390	),
	Cin=> Carry( 	2490	),
	Cout=> Carry( 	2491	),
	S=> E(	2452	));
			
  U2492	: Soma_AMA3_1 PORT MAP(
	A=> C(	2556	),
	B=>E(	2391	),
	Cin=> Carry( 	2491	),
	Cout=> Carry( 	2492	),
	S=> E(	2453	));
			
  U2493	: Soma_AMA3_1 PORT MAP(
	A=> C(	2557	),
	B=>E(	2392	),
	Cin=> Carry( 	2492	),
	Cout=> Carry( 	2493	),
	S=> E(	2454	));
			
  U2494	: Soma_AMA3_1 PORT MAP(
	A=> C(	2558	),
	B=>E(	2393	),
	Cin=> Carry( 	2493	),
	Cout=> Carry( 	2494	),
	S=> E(	2455	));
			
  U2495	: Soma_AMA3_1 PORT MAP(
	A=> C(	2559	),
	B=>Carry(	2431	),
	Cin=> Carry( 	2494	),
	Cout=> Carry( 	2495	),
	S=> E(	2456	));

			
  U2496	: Soma_AMA3_1 PORT MAP(
	A=> C(	2560	),
	B=>E(	2394	),
	Cin=> '0',
	Cout=> Carry( 	2496	),
	S=> R(	40	));
			
  U2497	: Soma_AMA3_1 PORT MAP(
	A=> C(	2561	),
	B=>E(	2395	),
	Cin=> Carry( 	2496	),
	Cout=> Carry( 	2497	),
	S=> E(	2457	));
			
  U2498	: Soma_AMA3_1 PORT MAP(
	A=> C(	2562	),
	B=>E(	2396	),
	Cin=> Carry( 	2497	),
	Cout=> Carry( 	2498	),
	S=> E(	2458	));
			
  U2499	: Soma_AMA3_1 PORT MAP(
	A=> C(	2563	),
	B=>E(	2397	),
	Cin=> Carry( 	2498	),
	Cout=> Carry( 	2499	),
	S=> E(	2459	));
			
  U2500	: Soma_AMA3_1 PORT MAP(
	A=> C(	2564	),
	B=>E(	2398	),
	Cin=> Carry( 	2499	),
	Cout=> Carry( 	2500	),
	S=> E(	2460	));
			
  U2501	: Soma_AMA3_1 PORT MAP(
	A=> C(	2565	),
	B=>E(	2399	),
	Cin=> Carry( 	2500	),
	Cout=> Carry( 	2501	),
	S=> E(	2461	));
			
  U2502	: Soma_AMA3_1 PORT MAP(
	A=> C(	2566	),
	B=>E(	2400	),
	Cin=> Carry( 	2501	),
	Cout=> Carry( 	2502	),
	S=> E(	2462	));
			
  U2503	: Soma_AMA3_1 PORT MAP(
	A=> C(	2567	),
	B=>E(	2401	),
	Cin=> Carry( 	2502	),
	Cout=> Carry( 	2503	),
	S=> E(	2463	));
			
  U2504	: Soma_AMA3_1 PORT MAP(
	A=> C(	2568	),
	B=>E(	2402	),
	Cin=> Carry( 	2503	),
	Cout=> Carry( 	2504	),
	S=> E(	2464	));
			
  U2505	: Soma_AMA3_1 PORT MAP(
	A=> C(	2569	),
	B=>E(	2403	),
	Cin=> Carry( 	2504	),
	Cout=> Carry( 	2505	),
	S=> E(	2465	));
			
  U2506	: Soma_AMA3_1 PORT MAP(
	A=> C(	2570	),
	B=>E(	2404	),
	Cin=> Carry( 	2505	),
	Cout=> Carry( 	2506	),
	S=> E(	2466	));
			
  U2507	: Soma_AMA3_1 PORT MAP(
	A=> C(	2571	),
	B=>E(	2405	),
	Cin=> Carry( 	2506	),
	Cout=> Carry( 	2507	),
	S=> E(	2467	));
			
  U2508	: Soma_AMA3_1 PORT MAP(
	A=> C(	2572	),
	B=>E(	2406	),
	Cin=> Carry( 	2507	),
	Cout=> Carry( 	2508	),
	S=> E(	2468	));
			
  U2509	: Soma_AMA3_1 PORT MAP(
	A=> C(	2573	),
	B=>E(	2407	),
	Cin=> Carry( 	2508	),
	Cout=> Carry( 	2509	),
	S=> E(	2469	));
			
  U2510	: Soma_AMA3_1 PORT MAP(
	A=> C(	2574	),
	B=>E(	2408	),
	Cin=> Carry( 	2509	),
	Cout=> Carry( 	2510	),
	S=> E(	2470	));
			
  U2511	: Soma_AMA3_1 PORT MAP(
	A=> C(	2575	),
	B=>E(	2409	),
	Cin=> Carry( 	2510	),
	Cout=> Carry( 	2511	),
	S=> E(	2471	));
			
  U2512	: Soma_AMA3_1 PORT MAP(
	A=> C(	2576	),
	B=>E(	2410	),
	Cin=> Carry( 	2511	),
	Cout=> Carry( 	2512	),
	S=> E(	2472	));
			
  U2513	: Soma_AMA3_1 PORT MAP(
	A=> C(	2577	),
	B=>E(	2411	),
	Cin=> Carry( 	2512	),
	Cout=> Carry( 	2513	),
	S=> E(	2473	));
			
  U2514	: Soma_AMA3_1 PORT MAP(
	A=> C(	2578	),
	B=>E(	2412	),
	Cin=> Carry( 	2513	),
	Cout=> Carry( 	2514	),
	S=> E(	2474	));
			
  U2515	: Soma_AMA3_1 PORT MAP(
	A=> C(	2579	),
	B=>E(	2413	),
	Cin=> Carry( 	2514	),
	Cout=> Carry( 	2515	),
	S=> E(	2475	));
			
  U2516	: Soma_AMA3_1 PORT MAP(
	A=> C(	2580	),
	B=>E(	2414	),
	Cin=> Carry( 	2515	),
	Cout=> Carry( 	2516	),
	S=> E(	2476	));
			
  U2517	: Soma_AMA3_1 PORT MAP(
	A=> C(	2581	),
	B=>E(	2415	),
	Cin=> Carry( 	2516	),
	Cout=> Carry( 	2517	),
	S=> E(	2477	));
			
  U2518	: Soma_AMA3_1 PORT MAP(
	A=> C(	2582	),
	B=>E(	2416	),
	Cin=> Carry( 	2517	),
	Cout=> Carry( 	2518	),
	S=> E(	2478	));
			
  U2519	: Soma_AMA3_1 PORT MAP(
	A=> C(	2583	),
	B=>E(	2417	),
	Cin=> Carry( 	2518	),
	Cout=> Carry( 	2519	),
	S=> E(	2479	));
			
  U2520	: Soma_AMA3_1 PORT MAP(
	A=> C(	2584	),
	B=>E(	2418	),
	Cin=> Carry( 	2519	),
	Cout=> Carry( 	2520	),
	S=> E(	2480	));
			
  U2521	: Soma_AMA3_1 PORT MAP(
	A=> C(	2585	),
	B=>E(	2419	),
	Cin=> Carry( 	2520	),
	Cout=> Carry( 	2521	),
	S=> E(	2481	));
			
  U2522	: Soma_AMA3_1 PORT MAP(
	A=> C(	2586	),
	B=>E(	2420	),
	Cin=> Carry( 	2521	),
	Cout=> Carry( 	2522	),
	S=> E(	2482	));
			
  U2523	: Soma_AMA3_1 PORT MAP(
	A=> C(	2587	),
	B=>E(	2421	),
	Cin=> Carry( 	2522	),
	Cout=> Carry( 	2523	),
	S=> E(	2483	));
			
  U2524	: Soma_AMA3_1 PORT MAP(
	A=> C(	2588	),
	B=>E(	2422	),
	Cin=> Carry( 	2523	),
	Cout=> Carry( 	2524	),
	S=> E(	2484	));
			
  U2525	: Soma_AMA3_1 PORT MAP(
	A=> C(	2589	),
	B=>E(	2423	),
	Cin=> Carry( 	2524	),
	Cout=> Carry( 	2525	),
	S=> E(	2485	));
			
  U2526	: Soma_AMA3_1 PORT MAP(
	A=> C(	2590	),
	B=>E(	2424	),
	Cin=> Carry( 	2525	),
	Cout=> Carry( 	2526	),
	S=> E(	2486	));
			
  U2527	: Soma_AMA3_1 PORT MAP(
	A=> C(	2591	),
	B=>E(	2425	),
	Cin=> Carry( 	2526	),
	Cout=> Carry( 	2527	),
	S=> E(	2487	));
			
  U2528	: Soma_AMA3_1 PORT MAP(
	A=> C(	2592	),
	B=>E(	2426	),
	Cin=> Carry( 	2527	),
	Cout=> Carry( 	2528	),
	S=> E(	2488	));
			
  U2529	: Soma_AMA3_1 PORT MAP(
	A=> C(	2593	),
	B=>E(	2427	),
	Cin=> Carry( 	2528	),
	Cout=> Carry( 	2529	),
	S=> E(	2489	));
			
  U2530	: Soma_AMA3_1 PORT MAP(
	A=> C(	2594	),
	B=>E(	2428	),
	Cin=> Carry( 	2529	),
	Cout=> Carry( 	2530	),
	S=> E(	2490	));
			
  U2531	: Soma_AMA3_1 PORT MAP(
	A=> C(	2595	),
	B=>E(	2429	),
	Cin=> Carry( 	2530	),
	Cout=> Carry( 	2531	),
	S=> E(	2491	));
			
  U2532	: Soma_AMA3_1 PORT MAP(
	A=> C(	2596	),
	B=>E(	2430	),
	Cin=> Carry( 	2531	),
	Cout=> Carry( 	2532	),
	S=> E(	2492	));
			
  U2533	: Soma_AMA3_1 PORT MAP(
	A=> C(	2597	),
	B=>E(	2431	),
	Cin=> Carry( 	2532	),
	Cout=> Carry( 	2533	),
	S=> E(	2493	));
			
  U2534	: Soma_AMA3_1 PORT MAP(
	A=> C(	2598	),
	B=>E(	2432	),
	Cin=> Carry( 	2533	),
	Cout=> Carry( 	2534	),
	S=> E(	2494	));
			
  U2535	: Soma_AMA3_1 PORT MAP(
	A=> C(	2599	),
	B=>E(	2433	),
	Cin=> Carry( 	2534	),
	Cout=> Carry( 	2535	),
	S=> E(	2495	));
			
  U2536	: Soma_AMA3_1 PORT MAP(
	A=> C(	2600	),
	B=>E(	2434	),
	Cin=> Carry( 	2535	),
	Cout=> Carry( 	2536	),
	S=> E(	2496	));
			
  U2537	: Soma_AMA3_1 PORT MAP(
	A=> C(	2601	),
	B=>E(	2435	),
	Cin=> Carry( 	2536	),
	Cout=> Carry( 	2537	),
	S=> E(	2497	));
			
  U2538	: Soma_AMA3_1 PORT MAP(
	A=> C(	2602	),
	B=>E(	2436	),
	Cin=> Carry( 	2537	),
	Cout=> Carry( 	2538	),
	S=> E(	2498	));
			
  U2539	: Soma_AMA3_1 PORT MAP(
	A=> C(	2603	),
	B=>E(	2437	),
	Cin=> Carry( 	2538	),
	Cout=> Carry( 	2539	),
	S=> E(	2499	));
			
  U2540	: Soma_AMA3_1 PORT MAP(
	A=> C(	2604	),
	B=>E(	2438	),
	Cin=> Carry( 	2539	),
	Cout=> Carry( 	2540	),
	S=> E(	2500	));
			
  U2541	: Soma_AMA3_1 PORT MAP(
	A=> C(	2605	),
	B=>E(	2439	),
	Cin=> Carry( 	2540	),
	Cout=> Carry( 	2541	),
	S=> E(	2501	));
			
  U2542	: Soma_AMA3_1 PORT MAP(
	A=> C(	2606	),
	B=>E(	2440	),
	Cin=> Carry( 	2541	),
	Cout=> Carry( 	2542	),
	S=> E(	2502	));
			
  U2543	: Soma_AMA3_1 PORT MAP(
	A=> C(	2607	),
	B=>E(	2441	),
	Cin=> Carry( 	2542	),
	Cout=> Carry( 	2543	),
	S=> E(	2503	));
			
  U2544	: Soma_AMA3_1 PORT MAP(
	A=> C(	2608	),
	B=>E(	2442	),
	Cin=> Carry( 	2543	),
	Cout=> Carry( 	2544	),
	S=> E(	2504	));
			
  U2545	: Soma_AMA3_1 PORT MAP(
	A=> C(	2609	),
	B=>E(	2443	),
	Cin=> Carry( 	2544	),
	Cout=> Carry( 	2545	),
	S=> E(	2505	));
			
  U2546	: Soma_AMA3_1 PORT MAP(
	A=> C(	2610	),
	B=>E(	2444	),
	Cin=> Carry( 	2545	),
	Cout=> Carry( 	2546	),
	S=> E(	2506	));
			
  U2547	: Soma_AMA3_1 PORT MAP(
	A=> C(	2611	),
	B=>E(	2445	),
	Cin=> Carry( 	2546	),
	Cout=> Carry( 	2547	),
	S=> E(	2507	));
			
  U2548	: Soma_AMA3_1 PORT MAP(
	A=> C(	2612	),
	B=>E(	2446	),
	Cin=> Carry( 	2547	),
	Cout=> Carry( 	2548	),
	S=> E(	2508	));
			
  U2549	: Soma_AMA3_1 PORT MAP(
	A=> C(	2613	),
	B=>E(	2447	),
	Cin=> Carry( 	2548	),
	Cout=> Carry( 	2549	),
	S=> E(	2509	));
			
  U2550	: Soma_AMA3_1 PORT MAP(
	A=> C(	2614	),
	B=>E(	2448	),
	Cin=> Carry( 	2549	),
	Cout=> Carry( 	2550	),
	S=> E(	2510	));
			
  U2551	: Soma_AMA3_1 PORT MAP(
	A=> C(	2615	),
	B=>E(	2449	),
	Cin=> Carry( 	2550	),
	Cout=> Carry( 	2551	),
	S=> E(	2511	));
			
  U2552	: Soma_AMA3_1 PORT MAP(
	A=> C(	2616	),
	B=>E(	2450	),
	Cin=> Carry( 	2551	),
	Cout=> Carry( 	2552	),
	S=> E(	2512	));
			
  U2553	: Soma_AMA3_1 PORT MAP(
	A=> C(	2617	),
	B=>E(	2451	),
	Cin=> Carry( 	2552	),
	Cout=> Carry( 	2553	),
	S=> E(	2513	));
			
  U2554	: Soma_AMA3_1 PORT MAP(
	A=> C(	2618	),
	B=>E(	2452	),
	Cin=> Carry( 	2553	),
	Cout=> Carry( 	2554	),
	S=> E(	2514	));
			
  U2555	: Soma_AMA3_1 PORT MAP(
	A=> C(	2619	),
	B=>E(	2453	),
	Cin=> Carry( 	2554	),
	Cout=> Carry( 	2555	),
	S=> E(	2515	));
			
  U2556	: Soma_AMA3_1 PORT MAP(
	A=> C(	2620	),
	B=>E(	2454	),
	Cin=> Carry( 	2555	),
	Cout=> Carry( 	2556	),
	S=> E(	2516	));
			
  U2557	: Soma_AMA3_1 PORT MAP(
	A=> C(	2621	),
	B=>E(	2455	),
	Cin=> Carry( 	2556	),
	Cout=> Carry( 	2557	),
	S=> E(	2517	));
			
  U2558	: Soma_AMA3_1 PORT MAP(
	A=> C(	2622	),
	B=>E(	2456	),
	Cin=> Carry( 	2557	),
	Cout=> Carry( 	2558	),
	S=> E(	2518	));
			
  U2559	: Soma_AMA3_1 PORT MAP(
	A => C(2623),
	B => Carry(2495),
	Cin => Carry(2558),
	Cout => Carry(2559),
	S => E(2519));

			
  U2560	: Soma_AMA3_1 PORT MAP(
	A=> C(	2624	),
	B=>E(	2457	),
	Cin=> '0'	,
	Cout=> Carry( 	2560	),
	S=> R(	41	));
			
  U2561	: Soma_AMA3_1 PORT MAP(
	A=> C(	2625	),
	B=>E(	2458	),
	Cin=> Carry( 	2560	),
	Cout=> Carry( 	2561	),
	S=> E(	2520	));
			
  U2562	: Soma_AMA3_1 PORT MAP(
	A=> C(	2626	),
	B=>E(	2459	),
	Cin=> Carry( 	2561	),
	Cout=> Carry( 	2562	),
	S=> E(	2521	));
			
  U2563	: Soma_AMA3_1 PORT MAP(
	A=> C(	2627	),
	B=>E(	2460	),
	Cin=> Carry( 	2562	),
	Cout=> Carry( 	2563	),
	S=> E(	2522	));
			
  U2564	: Soma_AMA3_1 PORT MAP(
	A=> C(	2628	),
	B=>E(	2461	),
	Cin=> Carry( 	2563	),
	Cout=> Carry( 	2564	),
	S=> E(	2523	));
			
  U2565	: Soma_AMA3_1 PORT MAP(
	A=> C(	2629	),
	B=>E(	2462	),
	Cin=> Carry( 	2564	),
	Cout=> Carry( 	2565	),
	S=> E(	2524	));
			
  U2566	: Soma_AMA3_1 PORT MAP(
	A=> C(	2630	),
	B=>E(	2463	),
	Cin=> Carry( 	2565	),
	Cout=> Carry( 	2566	),
	S=> E(	2525	));
			
  U2567	: Soma_AMA3_1 PORT MAP(
	A=> C(	2631	),
	B=>E(	2464	),
	Cin=> Carry( 	2566	),
	Cout=> Carry( 	2567	),
	S=> E(	2526	));
			
  U2568	: Soma_AMA3_1 PORT MAP(
	A=> C(	2632	),
	B=>E(	2465	),
	Cin=> Carry( 	2567	),
	Cout=> Carry( 	2568	),
	S=> E(	2527	));
			
  U2569	: Soma_AMA3_1 PORT MAP(
	A=> C(	2633	),
	B=>E(	2466	),
	Cin=> Carry( 	2568	),
	Cout=> Carry( 	2569	),
	S=> E(	2528	));
			
  U2570	: Soma_AMA3_1 PORT MAP(
	A=> C(	2634	),
	B=>E(	2467	),
	Cin=> Carry( 	2569	),
	Cout=> Carry( 	2570	),
	S=> E(	2529	));
			
  U2571	: Soma_AMA3_1 PORT MAP(
	A=> C(	2635	),
	B=>E(	2468	),
	Cin=> Carry( 	2570	),
	Cout=> Carry( 	2571	),
	S=> E(	2530	));
			
  U2572	: Soma_AMA3_1 PORT MAP(
	A=> C(	2636	),
	B=>E(	2469	),
	Cin=> Carry( 	2571	),
	Cout=> Carry( 	2572	),
	S=> E(	2531	));
			
  U2573	: Soma_AMA3_1 PORT MAP(
	A=> C(	2637	),
	B=>E(	2470	),
	Cin=> Carry( 	2572	),
	Cout=> Carry( 	2573	),
	S=> E(	2532	));
			
  U2574	: Soma_AMA3_1 PORT MAP(
	A=> C(	2638	),
	B=>E(	2471	),
	Cin=> Carry( 	2573	),
	Cout=> Carry( 	2574	),
	S=> E(	2533	));
			
  U2575	: Soma_AMA3_1 PORT MAP(
	A=> C(	2639	),
	B=>E(	2472	),
	Cin=> Carry( 	2574	),
	Cout=> Carry( 	2575	),
	S=> E(	2534	));
			
  U2576	: Soma_AMA3_1 PORT MAP(
	A=> C(	2640	),
	B=>E(	2473	),
	Cin=> Carry( 	2575	),
	Cout=> Carry( 	2576	),
	S=> E(	2535	));
			
  U2577	: Soma_AMA3_1 PORT MAP(
	A=> C(	2641	),
	B=>E(	2474	),
	Cin=> Carry( 	2576	),
	Cout=> Carry( 	2577	),
	S=> E(	2536	));
			
  U2578	: Soma_AMA3_1 PORT MAP(
	A=> C(	2642	),
	B=>E(	2475	),
	Cin=> Carry( 	2577	),
	Cout=> Carry( 	2578	),
	S=> E(	2537	));
			
  U2579	: Soma_AMA3_1 PORT MAP(
	A=> C(	2643	),
	B=>E(	2476	),
	Cin=> Carry( 	2578	),
	Cout=> Carry( 	2579	),
	S=> E(	2538	));
			
  U2580	: Soma_AMA3_1 PORT MAP(
	A=> C(	2644	),
	B=>E(	2477	),
	Cin=> Carry( 	2579	),
	Cout=> Carry( 	2580	),
	S=> E(	2539	));
			
  U2581	: Soma_AMA3_1 PORT MAP(
	A=> C(	2645	),
	B=>E(	2478	),
	Cin=> Carry( 	2580	),
	Cout=> Carry( 	2581	),
	S=> E(	2540	));
			
  U2582	: Soma_AMA3_1 PORT MAP(
	A=> C(	2646	),
	B=>E(	2479	),
	Cin=> Carry( 	2581	),
	Cout=> Carry( 	2582	),
	S=> E(	2541	));
			
  U2583	: Soma_AMA3_1 PORT MAP(
	A=> C(	2647	),
	B=>E(	2480	),
	Cin=> Carry( 	2582	),
	Cout=> Carry( 	2583	),
	S=> E(	2542	));
			
  U2584	: Soma_AMA3_1 PORT MAP(
	A=> C(	2648	),
	B=>E(	2481	),
	Cin=> Carry( 	2583	),
	Cout=> Carry( 	2584	),
	S=> E(	2543	));
			
  U2585	: Soma_AMA3_1 PORT MAP(
	A=> C(	2649	),
	B=>E(	2482	),
	Cin=> Carry( 	2584	),
	Cout=> Carry( 	2585	),
	S=> E(	2544	));
			
  U2586	: Soma_AMA3_1 PORT MAP(
	A=> C(	2650	),
	B=>E(	2483	),
	Cin=> Carry( 	2585	),
	Cout=> Carry( 	2586	),
	S=> E(	2545	));
			
  U2587	: Soma_AMA3_1 PORT MAP(
	A=> C(	2651	),
	B=>E(	2484	),
	Cin=> Carry( 	2586	),
	Cout=> Carry( 	2587	),
	S=> E(	2546	));
			
  U2588	: Soma_AMA3_1 PORT MAP(
	A=> C(	2652	),
	B=>E(	2485	),
	Cin=> Carry( 	2587	),
	Cout=> Carry( 	2588	),
	S=> E(	2547	));
			
  U2589	: Soma_AMA3_1 PORT MAP(
	A=> C(	2653	),
	B=>E(	2486	),
	Cin=> Carry( 	2588	),
	Cout=> Carry( 	2589	),
	S=> E(	2548	));
			
  U2590	: Soma_AMA3_1 PORT MAP(
	A=> C(	2654	),
	B=>E(	2487	),
	Cin=> Carry( 	2589	),
	Cout=> Carry( 	2590	),
	S=> E(	2549	));
			
  U2591	: Soma_AMA3_1 PORT MAP(
	A=> C(	2655	),
	B=>E(	2488	),
	Cin=> Carry( 	2590	),
	Cout=> Carry( 	2591	),
	S=> E(	2550	));
			
  U2592	: Soma_AMA3_1 PORT MAP(
	A=> C(	2656	),
	B=>E(	2489	),
	Cin=> Carry( 	2591	),
	Cout=> Carry( 	2592	),
	S=> E(	2551	));
			
  U2593	: Soma_AMA3_1 PORT MAP(
	A=> C(	2657	),
	B=>E(	2490	),
	Cin=> Carry( 	2592	),
	Cout=> Carry( 	2593	),
	S=> E(	2552	));
			
  U2594	: Soma_AMA3_1 PORT MAP(
	A=> C(	2658	),
	B=>E(	2491	),
	Cin=> Carry( 	2593	),
	Cout=> Carry( 	2594	),
	S=> E(	2553	));
			
  U2595	: Soma_AMA3_1 PORT MAP(
	A=> C(	2659	),
	B=>E(	2492	),
	Cin=> Carry( 	2594	),
	Cout=> Carry( 	2595	),
	S=> E(	2554	));
			
  U2596	: Soma_AMA3_1 PORT MAP(
	A=> C(	2660	),
	B=>E(	2493	),
	Cin=> Carry( 	2595	),
	Cout=> Carry( 	2596	),
	S=> E(	2555	));
			
  U2597	: Soma_AMA3_1 PORT MAP(
	A=> C(	2661	),
	B=>E(	2494	),
	Cin=> Carry( 	2596	),
	Cout=> Carry( 	2597	),
	S=> E(	2556	));
			
  U2598	: Soma_AMA3_1 PORT MAP(
	A=> C(	2662	),
	B=>E(	2495	),
	Cin=> Carry( 	2597	),
	Cout=> Carry( 	2598	),
	S=> E(	2557	));
			
  U2599	: Soma_AMA3_1 PORT MAP(
	A=> C(	2663	),
	B=>E(	2496	),
	Cin=> Carry( 	2598	),
	Cout=> Carry( 	2599	),
	S=> E(	2558	));
			
  U2600	: Soma_AMA3_1 PORT MAP(
	A=> C(	2664	),
	B=>E(	2497	),
	Cin=> Carry( 	2599	),
	Cout=> Carry( 	2600	),
	S=> E(	2559	));
			
  U2601	: Soma_AMA3_1 PORT MAP(
	A=> C(	2665	),
	B=>E(	2498	),
	Cin=> Carry( 	2600	),
	Cout=> Carry( 	2601	),
	S=> E(	2560	));
			
  U2602	: Soma_AMA3_1 PORT MAP(
	A=> C(	2666	),
	B=>E(	2499	),
	Cin=> Carry( 	2601	),
	Cout=> Carry( 	2602	),
	S=> E(	2561	));
			
  U2603	: Soma_AMA3_1 PORT MAP(
	A=> C(	2667	),
	B=>E(	2500	),
	Cin=> Carry( 	2602	),
	Cout=> Carry( 	2603	),
	S=> E(	2562	));
			
  U2604	: Soma_AMA3_1 PORT MAP(
	A=> C(	2668	),
	B=>E(	2501	),
	Cin=> Carry( 	2603	),
	Cout=> Carry( 	2604	),
	S=> E(	2563	));
			
  U2605	: Soma_AMA3_1 PORT MAP(
	A=> C(	2669	),
	B=>E(	2502	),
	Cin=> Carry( 	2604	),
	Cout=> Carry( 	2605	),
	S=> E(	2564	));
			
  U2606	: Soma_AMA3_1 PORT MAP(
	A=> C(	2670	),
	B=>E(	2503	),
	Cin=> Carry( 	2605	),
	Cout=> Carry( 	2606	),
	S=> E(	2565	));
			
  U2607	: Soma_AMA3_1 PORT MAP(
	A=> C(	2671	),
	B=>E(	2504	),
	Cin=> Carry( 	2606	),
	Cout=> Carry( 	2607	),
	S=> E(	2566	));
			
  U2608	: Soma_AMA3_1 PORT MAP(
	A=> C(	2672	),
	B=>E(	2505	),
	Cin=> Carry( 	2607	),
	Cout=> Carry( 	2608	),
	S=> E(	2567	));
			
  U2609	: Soma_AMA3_1 PORT MAP(
	A=> C(	2673	),
	B=>E(	2506	),
	Cin=> Carry( 	2608	),
	Cout=> Carry( 	2609	),
	S=> E(	2568	));
			
  U2610	: Soma_AMA3_1 PORT MAP(
	A=> C(	2674	),
	B=>E(	2507	),
	Cin=> Carry( 	2609	),
	Cout=> Carry( 	2610	),
	S=> E(	2569	));
			
  U2611	: Soma_AMA3_1 PORT MAP(
	A=> C(	2675	),
	B=>E(	2508	),
	Cin=> Carry( 	2610	),
	Cout=> Carry( 	2611	),
	S=> E(	2570	));
			
  U2612	: Soma_AMA3_1 PORT MAP(
	A=> C(	2676	),
	B=>E(	2509	),
	Cin=> Carry( 	2611	),
	Cout=> Carry( 	2612	),
	S=> E(	2571	));
			
  U2613	: Soma_AMA3_1 PORT MAP(
	A=> C(	2677	),
	B=>E(	2510	),
	Cin=> Carry( 	2612	),
	Cout=> Carry( 	2613	),
	S=> E(	2572	));
			
  U2614	: Soma_AMA3_1 PORT MAP(
	A=> C(	2678	),
	B=>E(	2511	),
	Cin=> Carry( 	2613	),
	Cout=> Carry( 	2614	),
	S=> E(	2573	));
			
  U2615	: Soma_AMA3_1 PORT MAP(
	A=> C(	2679	),
	B=>E(	2512	),
	Cin=> Carry( 	2614	),
	Cout=> Carry( 	2615	),
	S=> E(	2574	));
			
  U2616	: Soma_AMA3_1 PORT MAP(
	A=> C(	2680	),
	B=>E(	2513	),
	Cin=> Carry( 	2615	),
	Cout=> Carry( 	2616	),
	S=> E(	2575	));
			
  U2617	: Soma_AMA3_1 PORT MAP(
	A=> C(	2681	),
	B=>E(	2514	),
	Cin=> Carry( 	2616	),
	Cout=> Carry( 	2617	),
	S=> E(	2576	));
			
  U2618	: Soma_AMA3_1 PORT MAP(
	A=> C(	2682	),
	B=>E(	2515	),
	Cin=> Carry( 	2617	),
	Cout=> Carry( 	2618	),
	S=> E(	2577	));
			
  U2619	: Soma_AMA3_1 PORT MAP(
	A=> C(	2683	),
	B=>E(	2516	),
	Cin=> Carry( 	2618	),
	Cout=> Carry( 	2619	),
	S=> E(	2578	));
			
  U2620	: Soma_AMA3_1 PORT MAP(
	A=> C(	2684	),
	B=>E(	2517	),
	Cin=> Carry( 	2619	),
	Cout=> Carry( 	2620	),
	S=> E(	2579	));
			
  U2621	: Soma_AMA3_1 PORT MAP(
	A=> C(	2685	),
	B=>E(	2518	),
	Cin=> Carry( 	2620	),
	Cout=> Carry( 	2621	),
	S=> E(	2580	));
			
  U2622	: Soma_AMA3_1 PORT MAP(
	A=> C(	2686	),
	B=>E(	2519	),
	Cin=> Carry( 	2621	),
	Cout=> Carry( 	2622	),
	S=> E(	2581	));
			
  U2623	: Soma_AMA3_1 PORT MAP(
	A=> C(	2687	),
	B=>Carry(	2559	),
	Cin=> Carry( 	2622	),
	Cout=> Carry( 	2623	),
	S=> E(	2582	));

			
  U2624	: Soma_AMA3_1 PORT MAP(
	A=> C(	2688	),
	B=>E(	2520	),
	Cin=> '0'	,
	Cout=> Carry( 	2624	),
	S=> R(	42	));
			
  U2625	: Soma_AMA3_1 PORT MAP(
	A=> C(	2689	),
	B=>E(	2521	),
	Cin=> Carry( 	2624	),
	Cout=> Carry( 	2625	),
	S=> E(	2583	));
			
  U2626	: Soma_AMA3_1 PORT MAP(
	A=> C(	2690	),
	B=>E(	2522	),
	Cin=> Carry( 	2625	),
	Cout=> Carry( 	2626	),
	S=> E(	2584	));
			
  U2627	: Soma_AMA3_1 PORT MAP(
	A=> C(	2691	),
	B=>E(	2523	),
	Cin=> Carry( 	2626	),
	Cout=> Carry( 	2627	),
	S=> E(	2585	));
			
  U2628	: Soma_AMA3_1 PORT MAP(
	A=> C(	2692	),
	B=>E(	2524	),
	Cin=> Carry( 	2627	),
	Cout=> Carry( 	2628	),
	S=> E(	2586	));
			
  U2629	: Soma_AMA3_1 PORT MAP(
	A=> C(	2693	),
	B=>E(	2525	),
	Cin=> Carry( 	2628	),
	Cout=> Carry( 	2629	),
	S=> E(	2587	));
			
  U2630	: Soma_AMA3_1 PORT MAP(
	A=> C(	2694	),
	B=>E(	2526	),
	Cin=> Carry( 	2629	),
	Cout=> Carry( 	2630	),
	S=> E(	2588	));
			
  U2631	: Soma_AMA3_1 PORT MAP(
	A=> C(	2695	),
	B=>E(	2527	),
	Cin=> Carry( 	2630	),
	Cout=> Carry( 	2631	),
	S=> E(	2589	));
			
  U2632	: Soma_AMA3_1 PORT MAP(
	A=> C(	2696	),
	B=>E(	2528	),
	Cin=> Carry( 	2631	),
	Cout=> Carry( 	2632	),
	S=> E(	2590	));
			
  U2633	: Soma_AMA3_1 PORT MAP(
	A=> C(	2697	),
	B=>E(	2529	),
	Cin=> Carry( 	2632	),
	Cout=> Carry( 	2633	),
	S=> E(	2591	));
			
  U2634	: Soma_AMA3_1 PORT MAP(
	A=> C(	2698	),
	B=>E(	2530	),
	Cin=> Carry( 	2633	),
	Cout=> Carry( 	2634	),
	S=> E(	2592	));
			
  U2635	: Soma_AMA3_1 PORT MAP(
	A=> C(	2699	),
	B=>E(	2531	),
	Cin=> Carry( 	2634	),
	Cout=> Carry( 	2635	),
	S=> E(	2593	));
			
  U2636	: Soma_AMA3_1 PORT MAP(
	A=> C(	2700	),
	B=>E(	2532	),
	Cin=> Carry( 	2635	),
	Cout=> Carry( 	2636	),
	S=> E(	2594	));
			
  U2637	: Soma_AMA3_1 PORT MAP(
	A=> C(	2701	),
	B=>E(	2533	),
	Cin=> Carry( 	2636	),
	Cout=> Carry( 	2637	),
	S=> E(	2595	));
			
  U2638	: Soma_AMA3_1 PORT MAP(
	A=> C(	2702	),
	B=>E(	2534	),
	Cin=> Carry( 	2637	),
	Cout=> Carry( 	2638	),
	S=> E(	2596	));
			
  U2639	: Soma_AMA3_1 PORT MAP(
	A=> C(	2703	),
	B=>E(	2535	),
	Cin=> Carry( 	2638	),
	Cout=> Carry( 	2639	),
	S=> E(	2597	));
			
  U2640	: Soma_AMA3_1 PORT MAP(
	A=> C(	2704	),
	B=>E(	2536	),
	Cin=> Carry( 	2639	),
	Cout=> Carry( 	2640	),
	S=> E(	2598	));
			
  U2641	: Soma_AMA3_1 PORT MAP(
	A=> C(	2705	),
	B=>E(	2537	),
	Cin=> Carry( 	2640	),
	Cout=> Carry( 	2641	),
	S=> E(	2599	));
			
  U2642	: Soma_AMA3_1 PORT MAP(
	A=> C(	2706	),
	B=>E(	2538	),
	Cin=> Carry( 	2641	),
	Cout=> Carry( 	2642	),
	S=> E(	2600	));
			
  U2643	: Soma_AMA3_1 PORT MAP(
	A=> C(	2707	),
	B=>E(	2539	),
	Cin=> Carry( 	2642	),
	Cout=> Carry( 	2643	),
	S=> E(	2601	));
			
  U2644	: Soma_AMA3_1 PORT MAP(
	A=> C(	2708	),
	B=>E(	2540	),
	Cin=> Carry( 	2643	),
	Cout=> Carry( 	2644	),
	S=> E(	2602	));
			
  U2645	: Soma_AMA3_1 PORT MAP(
	A=> C(	2709	),
	B=>E(	2541	),
	Cin=> Carry( 	2644	),
	Cout=> Carry( 	2645	),
	S=> E(	2603	));
			
  U2646	: Soma_AMA3_1 PORT MAP(
	A=> C(	2710	),
	B=>E(	2542	),
	Cin=> Carry( 	2645	),
	Cout=> Carry( 	2646	),
	S=> E(	2604	));
			
  U2647	: Soma_AMA3_1 PORT MAP(
	A=> C(	2711	),
	B=>E(	2543	),
	Cin=> Carry( 	2646	),
	Cout=> Carry( 	2647	),
	S=> E(	2605	));
			
  U2648	: Soma_AMA3_1 PORT MAP(
	A=> C(	2712	),
	B=>E(	2544	),
	Cin=> Carry( 	2647	),
	Cout=> Carry( 	2648	),
	S=> E(	2606	));
			
  U2649	: Soma_AMA3_1 PORT MAP(
	A=> C(	2713	),
	B=>E(	2545	),
	Cin=> Carry( 	2648	),
	Cout=> Carry( 	2649	),
	S=> E(	2607	));
			
  U2650	: Soma_AMA3_1 PORT MAP(
	A=> C(	2714	),
	B=>E(	2546	),
	Cin=> Carry( 	2649	),
	Cout=> Carry( 	2650	),
	S=> E(	2608	));
			
  U2651	: Soma_AMA3_1 PORT MAP(
	A=> C(	2715	),
	B=>E(	2547	),
	Cin=> Carry( 	2650	),
	Cout=> Carry( 	2651	),
	S=> E(	2609	));
			
  U2652	: Soma_AMA3_1 PORT MAP(
	A=> C(	2716	),
	B=>E(	2548	),
	Cin=> Carry( 	2651	),
	Cout=> Carry( 	2652	),
	S=> E(	2610	));
			
  U2653	: Soma_AMA3_1 PORT MAP(
	A=> C(	2717	),
	B=>E(	2549	),
	Cin=> Carry( 	2652	),
	Cout=> Carry( 	2653	),
	S=> E(	2611	));
			
  U2654	: Soma_AMA3_1 PORT MAP(
	A=> C(	2718	),
	B=>E(	2550	),
	Cin=> Carry( 	2653	),
	Cout=> Carry( 	2654	),
	S=> E(	2612	));
			
  U2655	: Soma_AMA3_1 PORT MAP(
	A=> C(	2719	),
	B=>E(	2551	),
	Cin=> Carry( 	2654	),
	Cout=> Carry( 	2655	),
	S=> E(	2613	));
			
  U2656	: Soma_AMA3_1 PORT MAP(
	A=> C(	2720	),
	B=>E(	2552	),
	Cin=> Carry( 	2655	),
	Cout=> Carry( 	2656	),
	S=> E(	2614	));
			
  U2657	: Soma_AMA3_1 PORT MAP(
	A=> C(	2721	),
	B=>E(	2553	),
	Cin=> Carry( 	2656	),
	Cout=> Carry( 	2657	),
	S=> E(	2615	));
			
  U2658	: Soma_AMA3_1 PORT MAP(
	A=> C(	2722	),
	B=>E(	2554	),
	Cin=> Carry( 	2657	),
	Cout=> Carry( 	2658	),
	S=> E(	2616	));
			
  U2659	: Soma_AMA3_1 PORT MAP(
	A=> C(	2723	),
	B=>E(	2555	),
	Cin=> Carry( 	2658	),
	Cout=> Carry( 	2659	),
	S=> E(	2617	));
			
  U2660	: Soma_AMA3_1 PORT MAP(
	A=> C(	2724	),
	B=>E(	2556	),
	Cin=> Carry( 	2659	),
	Cout=> Carry( 	2660	),
	S=> E(	2618	));
			
  U2661	: Soma_AMA3_1 PORT MAP(
	A=> C(	2725	),
	B=>E(	2557	),
	Cin=> Carry( 	2660	),
	Cout=> Carry( 	2661	),
	S=> E(	2619	));
			
  U2662	: Soma_AMA3_1 PORT MAP(
	A=> C(	2726	),
	B=>E(	2558	),
	Cin=> Carry( 	2661	),
	Cout=> Carry( 	2662	),
	S=> E(	2620	));
			
  U2663	: Soma_AMA3_1 PORT MAP(
	A=> C(	2727	),
	B=>E(	2559	),
	Cin=> Carry( 	2662	),
	Cout=> Carry( 	2663	),
	S=> E(	2621	));
			
  U2664	: Soma_AMA3_1 PORT MAP(
	A=> C(	2728	),
	B=>E(	2560	),
	Cin=> Carry( 	2663	),
	Cout=> Carry( 	2664	),
	S=> E(	2622	));
			
  U2665	: Soma_AMA3_1 PORT MAP(
	A=> C(	2729	),
	B=>E(	2561	),
	Cin=> Carry( 	2664	),
	Cout=> Carry( 	2665	),
	S=> E(	2623	));
			
  U2666	: Soma_AMA3_1 PORT MAP(
	A=> C(	2730	),
	B=>E(	2562	),
	Cin=> Carry( 	2665	),
	Cout=> Carry( 	2666	),
	S=> E(	2624	));
			
  U2667	: Soma_AMA3_1 PORT MAP(
	A=> C(	2731	),
	B=>E(	2563	),
	Cin=> Carry( 	2666	),
	Cout=> Carry( 	2667	),
	S=> E(	2625	));
			
  U2668	: Soma_AMA3_1 PORT MAP(
	A=> C(	2732	),
	B=>E(	2564	),
	Cin=> Carry( 	2667	),
	Cout=> Carry( 	2668	),
	S=> E(	2626	));
			
  U2669	: Soma_AMA3_1 PORT MAP(
	A=> C(	2733	),
	B=>E(	2565	),
	Cin=> Carry( 	2668	),
	Cout=> Carry( 	2669	),
	S=> E(	2627	));
			
  U2670	: Soma_AMA3_1 PORT MAP(
	A=> C(	2734	),
	B=>E(	2566	),
	Cin=> Carry( 	2669	),
	Cout=> Carry( 	2670	),
	S=> E(	2628	));
			
  U2671	: Soma_AMA3_1 PORT MAP(
	A=> C(	2735	),
	B=>E(	2567	),
	Cin=> Carry( 	2670	),
	Cout=> Carry( 	2671	),
	S=> E(	2629	));
			
  U2672	: Soma_AMA3_1 PORT MAP(
	A=> C(	2736	),
	B=>E(	2568	),
	Cin=> Carry( 	2671	),
	Cout=> Carry( 	2672	),
	S=> E(	2630	));
			
  U2673	: Soma_AMA3_1 PORT MAP(
	A=> C(	2737	),
	B=>E(	2569	),
	Cin=> Carry( 	2672	),
	Cout=> Carry( 	2673	),
	S=> E(	2631	));
			
  U2674	: Soma_AMA3_1 PORT MAP(
	A=> C(	2738	),
	B=>E(	2570	),
	Cin=> Carry( 	2673	),
	Cout=> Carry( 	2674	),
	S=> E(	2632	));
			
  U2675	: Soma_AMA3_1 PORT MAP(
	A=> C(	2739	),
	B=>E(	2571	),
	Cin=> Carry( 	2674	),
	Cout=> Carry( 	2675	),
	S=> E(	2633	));
			
  U2676	: Soma_AMA3_1 PORT MAP(
	A=> C(	2740	),
	B=>E(	2572	),
	Cin=> Carry( 	2675	),
	Cout=> Carry( 	2676	),
	S=> E(	2634	));
			
  U2677	: Soma_AMA3_1 PORT MAP(
	A=> C(	2741	),
	B=>E(	2573	),
	Cin=> Carry( 	2676	),
	Cout=> Carry( 	2677	),
	S=> E(	2635	));
			
  U2678	: Soma_AMA3_1 PORT MAP(
	A=> C(	2742	),
	B=>E(	2574	),
	Cin=> Carry( 	2677	),
	Cout=> Carry( 	2678	),
	S=> E(	2636	));
			
  U2679	: Soma_AMA3_1 PORT MAP(
	A=> C(	2743	),
	B=>E(	2575	),
	Cin=> Carry( 	2678	),
	Cout=> Carry( 	2679	),
	S=> E(	2637	));
			
  U2680	: Soma_AMA3_1 PORT MAP(
	A=> C(	2744	),
	B=>E(	2576	),
	Cin=> Carry( 	2679	),
	Cout=> Carry( 	2680	),
	S=> E(	2638	));
			
  U2681	: Soma_AMA3_1 PORT MAP(
	A=> C(	2745	),
	B=>E(	2577	),
	Cin=> Carry( 	2680	),
	Cout=> Carry( 	2681	),
	S=> E(	2639	));
			
  U2682	: Soma_AMA3_1 PORT MAP(
	A=> C(	2746	),
	B=>E(	2578	),
	Cin=> Carry( 	2681	),
	Cout=> Carry( 	2682	),
	S=> E(	2640	));
			
  U2683	: Soma_AMA3_1 PORT MAP(
	A=> C(	2747	),
	B=>E(	2579	),
	Cin=> Carry( 	2682	),
	Cout=> Carry( 	2683	),
	S=> E(	2641	));
			
  U2684	: Soma_AMA3_1 PORT MAP(
	A=> C(	2748	),
	B=>E(	2580	),
	Cin=> Carry( 	2683	),
	Cout=> Carry( 	2684	),
	S=> E(	2642	));
			
  U2685	: Soma_AMA3_1 PORT MAP(
	A=> C(	2749	),
	B=>E(	2581	),
	Cin=> Carry( 	2684	),
	Cout=> Carry( 	2685	),
	S=> E(	2643	));
			
  U2686	: Soma_AMA3_1 PORT MAP(
	A=> C(	2750	),
	B=>E(	2582	),
	Cin=> Carry( 	2685	),
	Cout=> Carry( 	2686	),
	S=> E(	2644	));
			
  U2687	: Soma_AMA3_1 PORT MAP(
	A=> C(	2751	),
	B=>Carry(	2623	),
	Cin=> Carry( 	2686	),
	Cout=> Carry( 	2687	),
	S=> E(	2645	));

			
  U2688	: Soma_AMA3_1 PORT MAP(
	A=> C(	2752	),
	B=>E(	2583	),
	Cin=> '0',
	Cout=> Carry( 	2688	),
	S=> R(	43	));
			
  U2689	: Soma_AMA3_1 PORT MAP(
	A=> C(	2753	),
	B=>E(	2584	),
	Cin=> Carry( 	2688	),
	Cout=> Carry( 	2689	),
	S=> E(	2646	));
			
  U2690	: Soma_AMA3_1 PORT MAP(
	A=> C(	2754	),
	B=>E(	2585	),
	Cin=> Carry( 	2689	),
	Cout=> Carry( 	2690	),
	S=> E(	2647	));
			
  U2691	: Soma_AMA3_1 PORT MAP(
	A=> C(	2755	),
	B=>E(	2586	),
	Cin=> Carry( 	2690	),
	Cout=> Carry( 	2691	),
	S=> E(	2648	));
			
  U2692	: Soma_AMA3_1 PORT MAP(
	A=> C(	2756	),
	B=>E(	2587	),
	Cin=> Carry( 	2691	),
	Cout=> Carry( 	2692	),
	S=> E(	2649	));
			
  U2693	: Soma_AMA3_1 PORT MAP(
	A=> C(	2757	),
	B=>E(	2588	),
	Cin=> Carry( 	2692	),
	Cout=> Carry( 	2693	),
	S=> E(	2650	));
			
  U2694	: Soma_AMA3_1 PORT MAP(
	A=> C(	2758	),
	B=>E(	2589	),
	Cin=> Carry( 	2693	),
	Cout=> Carry( 	2694	),
	S=> E(	2651	));
			
  U2695	: Soma_AMA3_1 PORT MAP(
	A=> C(	2759	),
	B=>E(	2590	),
	Cin=> Carry( 	2694	),
	Cout=> Carry( 	2695	),
	S=> E(	2652	));
			
  U2696	: Soma_AMA3_1 PORT MAP(
	A=> C(	2760	),
	B=>E(	2591	),
	Cin=> Carry( 	2695	),
	Cout=> Carry( 	2696	),
	S=> E(	2653	));
			
  U2697	: Soma_AMA3_1 PORT MAP(
	A=> C(	2761	),
	B=>E(	2592	),
	Cin=> Carry( 	2696	),
	Cout=> Carry( 	2697	),
	S=> E(	2654	));
			
  U2698	: Soma_AMA3_1 PORT MAP(
	A=> C(	2762	),
	B=>E(	2593	),
	Cin=> Carry( 	2697	),
	Cout=> Carry( 	2698	),
	S=> E(	2655	));
			
  U2699	: Soma_AMA3_1 PORT MAP(
	A=> C(	2763	),
	B=>E(	2594	),
	Cin=> Carry( 	2698	),
	Cout=> Carry( 	2699	),
	S=> E(	2656	));
			
  U2700	: Soma_AMA3_1 PORT MAP(
	A=> C(	2764	),
	B=>E(	2595	),
	Cin=> Carry( 	2699	),
	Cout=> Carry( 	2700	),
	S=> E(	2657	));
			
  U2701	: Soma_AMA3_1 PORT MAP(
	A=> C(	2765	),
	B=>E(	2596	),
	Cin=> Carry( 	2700	),
	Cout=> Carry( 	2701	),
	S=> E(	2658	));
			
  U2702	: Soma_AMA3_1 PORT MAP(
	A=> C(	2766	),
	B=>E(	2597	),
	Cin=> Carry( 	2701	),
	Cout=> Carry( 	2702	),
	S=> E(	2659	));
			
  U2703	: Soma_AMA3_1 PORT MAP(
	A=> C(	2767	),
	B=>E(	2598	),
	Cin=> Carry( 	2702	),
	Cout=> Carry( 	2703	),
	S=> E(	2660	));
			
  U2704	: Soma_AMA3_1 PORT MAP(
	A=> C(	2768	),
	B=>E(	2599	),
	Cin=> Carry( 	2703	),
	Cout=> Carry( 	2704	),
	S=> E(	2661	));
			
  U2705	: Soma_AMA3_1 PORT MAP(
	A=> C(	2769	),
	B=>E(	2600	),
	Cin=> Carry( 	2704	),
	Cout=> Carry( 	2705	),
	S=> E(	2662	));
			
  U2706	: Soma_AMA3_1 PORT MAP(
	A=> C(	2770	),
	B=>E(	2601	),
	Cin=> Carry( 	2705	),
	Cout=> Carry( 	2706	),
	S=> E(	2663	));
			
  U2707	: Soma_AMA3_1 PORT MAP(
	A=> C(	2771	),
	B=>E(	2602	),
	Cin=> Carry( 	2706	),
	Cout=> Carry( 	2707	),
	S=> E(	2664	));
			
  U2708	: Soma_AMA3_1 PORT MAP(
	A=> C(	2772	),
	B=>E(	2603	),
	Cin=> Carry( 	2707	),
	Cout=> Carry( 	2708	),
	S=> E(	2665	));
			
  U2709	: Soma_AMA3_1 PORT MAP(
	A=> C(	2773	),
	B=>E(	2604	),
	Cin=> Carry( 	2708	),
	Cout=> Carry( 	2709	),
	S=> E(	2666	));
			
  U2710	: Soma_AMA3_1 PORT MAP(
	A=> C(	2774	),
	B=>E(	2605	),
	Cin=> Carry( 	2709	),
	Cout=> Carry( 	2710	),
	S=> E(	2667	));
			
  U2711	: Soma_AMA3_1 PORT MAP(
	A=> C(	2775	),
	B=>E(	2606	),
	Cin=> Carry( 	2710	),
	Cout=> Carry( 	2711	),
	S=> E(	2668	));
			
  U2712	: Soma_AMA3_1 PORT MAP(
	A=> C(	2776	),
	B=>E(	2607	),
	Cin=> Carry( 	2711	),
	Cout=> Carry( 	2712	),
	S=> E(	2669	));
			
  U2713	: Soma_AMA3_1 PORT MAP(
	A=> C(	2777	),
	B=>E(	2608	),
	Cin=> Carry( 	2712	),
	Cout=> Carry( 	2713	),
	S=> E(	2670	));
			
  U2714	: Soma_AMA3_1 PORT MAP(
	A=> C(	2778	),
	B=>E(	2609	),
	Cin=> Carry( 	2713	),
	Cout=> Carry( 	2714	),
	S=> E(	2671	));
			
  U2715	: Soma_AMA3_1 PORT MAP(
	A=> C(	2779	),
	B=>E(	2610	),
	Cin=> Carry( 	2714	),
	Cout=> Carry( 	2715	),
	S=> E(	2672	));
			
  U2716	: Soma_AMA3_1 PORT MAP(
	A=> C(	2780	),
	B=>E(	2611	),
	Cin=> Carry( 	2715	),
	Cout=> Carry( 	2716	),
	S=> E(	2673	));
			
  U2717	: Soma_AMA3_1 PORT MAP(
	A=> C(	2781	),
	B=>E(	2612	),
	Cin=> Carry( 	2716	),
	Cout=> Carry( 	2717	),
	S=> E(	2674	));
			
  U2718	: Soma_AMA3_1 PORT MAP(
	A=> C(	2782	),
	B=>E(	2613	),
	Cin=> Carry( 	2717	),
	Cout=> Carry( 	2718	),
	S=> E(	2675	));
			
  U2719	: Soma_AMA3_1 PORT MAP(
	A=> C(	2783	),
	B=>E(	2614	),
	Cin=> Carry( 	2718	),
	Cout=> Carry( 	2719	),
	S=> E(	2676	));
			
  U2720	: Soma_AMA3_1 PORT MAP(
	A=> C(	2784	),
	B=>E(	2615	),
	Cin=> Carry( 	2719	),
	Cout=> Carry( 	2720	),
	S=> E(	2677	));
			
  U2721	: Soma_AMA3_1 PORT MAP(
	A=> C(	2785	),
	B=>E(	2616	),
	Cin=> Carry( 	2720	),
	Cout=> Carry( 	2721	),
	S=> E(	2678	));
			
  U2722	: Soma_AMA3_1 PORT MAP(
	A=> C(	2786	),
	B=>E(	2617	),
	Cin=> Carry( 	2721	),
	Cout=> Carry( 	2722	),
	S=> E(	2679	));
			
  U2723	: Soma_AMA3_1 PORT MAP(
	A=> C(	2787	),
	B=>E(	2618	),
	Cin=> Carry( 	2722	),
	Cout=> Carry( 	2723	),
	S=> E(	2680	));
			
  U2724	: Soma_AMA3_1 PORT MAP(
	A=> C(	2788	),
	B=>E(	2619	),
	Cin=> Carry( 	2723	),
	Cout=> Carry( 	2724	),
	S=> E(	2681	));
			
  U2725	: Soma_AMA3_1 PORT MAP(
	A=> C(	2789	),
	B=>E(	2620	),
	Cin=> Carry( 	2724	),
	Cout=> Carry( 	2725	),
	S=> E(	2682	));
			
  U2726	: Soma_AMA3_1 PORT MAP(
	A=> C(	2790	),
	B=>E(	2621	),
	Cin=> Carry( 	2725	),
	Cout=> Carry( 	2726	),
	S=> E(	2683	));
			
  U2727	: Soma_AMA3_1 PORT MAP(
	A=> C(	2791	),
	B=>E(	2622	),
	Cin=> Carry( 	2726	),
	Cout=> Carry( 	2727	),
	S=> E(	2684	));
			
  U2728	: Soma_AMA3_1 PORT MAP(
	A=> C(	2792	),
	B=>E(	2623	),
	Cin=> Carry( 	2727	),
	Cout=> Carry( 	2728	),
	S=> E(	2685	));
			
  U2729	: Soma_AMA3_1 PORT MAP(
	A=> C(	2793	),
	B=>E(	2624	),
	Cin=> Carry( 	2728	),
	Cout=> Carry( 	2729	),
	S=> E(	2686	));
			
  U2730	: Soma_AMA3_1 PORT MAP(
	A=> C(	2794	),
	B=>E(	2625	),
	Cin=> Carry( 	2729	),
	Cout=> Carry( 	2730	),
	S=> E(	2687	));
			
  U2731	: Soma_AMA3_1 PORT MAP(
	A=> C(	2795	),
	B=>E(	2626	),
	Cin=> Carry( 	2730	),
	Cout=> Carry( 	2731	),
	S=> E(	2688	));
			
  U2732	: Soma_AMA3_1 PORT MAP(
	A=> C(	2796	),
	B=>E(	2627	),
	Cin=> Carry( 	2731	),
	Cout=> Carry( 	2732	),
	S=> E(	2689	));
			
  U2733	: Soma_AMA3_1 PORT MAP(
	A=> C(	2797	),
	B=>E(	2628	),
	Cin=> Carry( 	2732	),
	Cout=> Carry( 	2733	),
	S=> E(	2690	));
			
  U2734	: Soma_AMA3_1 PORT MAP(
	A=> C(	2798	),
	B=>E(	2629	),
	Cin=> Carry( 	2733	),
	Cout=> Carry( 	2734	),
	S=> E(	2691	));
			
  U2735	: Soma_AMA3_1 PORT MAP(
	A=> C(	2799	),
	B=>E(	2630	),
	Cin=> Carry( 	2734	),
	Cout=> Carry( 	2735	),
	S=> E(	2692	));
			
  U2736	: Soma_AMA3_1 PORT MAP(
	A=> C(	2800	),
	B=>E(	2631	),
	Cin=> Carry( 	2735	),
	Cout=> Carry( 	2736	),
	S=> E(	2693	));
			
  U2737	: Soma_AMA3_1 PORT MAP(
	A=> C(	2801	),
	B=>E(	2632	),
	Cin=> Carry( 	2736	),
	Cout=> Carry( 	2737	),
	S=> E(	2694	));
			
  U2738	: Soma_AMA3_1 PORT MAP(
	A=> C(	2802	),
	B=>E(	2633	),
	Cin=> Carry( 	2737	),
	Cout=> Carry( 	2738	),
	S=> E(	2695	));
			
  U2739	: Soma_AMA3_1 PORT MAP(
	A=> C(	2803	),
	B=>E(	2634	),
	Cin=> Carry( 	2738	),
	Cout=> Carry( 	2739	),
	S=> E(	2696	));
			
  U2740	: Soma_AMA3_1 PORT MAP(
	A=> C(	2804	),
	B=>E(	2635	),
	Cin=> Carry( 	2739	),
	Cout=> Carry( 	2740	),
	S=> E(	2697	));
			
  U2741	: Soma_AMA3_1 PORT MAP(
	A=> C(	2805	),
	B=>E(	2636	),
	Cin=> Carry( 	2740	),
	Cout=> Carry( 	2741	),
	S=> E(	2698	));
			
  U2742	: Soma_AMA3_1 PORT MAP(
	A=> C(	2806	),
	B=>E(	2637	),
	Cin=> Carry( 	2741	),
	Cout=> Carry( 	2742	),
	S=> E(	2699	));
			
  U2743	: Soma_AMA3_1 PORT MAP(
	A=> C(	2807	),
	B=>E(	2638	),
	Cin=> Carry( 	2742	),
	Cout=> Carry( 	2743	),
	S=> E(	2700	));
			
  U2744	: Soma_AMA3_1 PORT MAP(
	A=> C(	2808	),
	B=>E(	2639	),
	Cin=> Carry( 	2743	),
	Cout=> Carry( 	2744	),
	S=> E(	2701	));
			
  U2745	: Soma_AMA3_1 PORT MAP(
	A=> C(	2809	),
	B=>E(	2640	),
	Cin=> Carry( 	2744	),
	Cout=> Carry( 	2745	),
	S=> E(	2702	));
			
  U2746	: Soma_AMA3_1 PORT MAP(
	A=> C(	2810	),
	B=>E(	2641	),
	Cin=> Carry( 	2745	),
	Cout=> Carry( 	2746	),
	S=> E(	2703	));
			
  U2747	: Soma_AMA3_1 PORT MAP(
	A=> C(	2811	),
	B=>E(	2642	),
	Cin=> Carry( 	2746	),
	Cout=> Carry( 	2747	),
	S=> E(	2704	));
			
  U2748	: Soma_AMA3_1 PORT MAP(
	A=> C(	2812	),
	B=>E(	2643	),
	Cin=> Carry( 	2747	),
	Cout=> Carry( 	2748	),
	S=> E(	2705	));
			
  U2749	: Soma_AMA3_1 PORT MAP(
	A=> C(	2813	),
	B=>E(	2644	),
	Cin=> Carry( 	2748	),
	Cout=> Carry( 	2749	),
	S=> E(	2706	));
			
  U2750	: Soma_AMA3_1 PORT MAP(
	A=> C(	2814	),
	B=>E(	2645	),
	Cin=> Carry( 	2749	),
	Cout=> Carry( 	2750	),
	S=> E(	2707	));
			
  U2751	: Soma_AMA3_1 PORT MAP(
	A=> C(	2815	),
	B=>Carry(	2687	),
	Cin=> Carry( 	2750	),
	Cout=> Carry( 	2751	),
	S=> E(	2708	));

			
  U2752	: Soma_AMA3_1 PORT MAP(
	A=> C(	2816	),
	B=>E(	2646	),
	Cin=> '0'	,
	Cout=> Carry( 	2752	),
	S=> R(	44	));
			
  U2753	: Soma_AMA3_1 PORT MAP(
	A=> C(	2817	),
	B=>E(	2647	),
	Cin=> Carry( 	2752	),
	Cout=> Carry( 	2753	),
	S=> E(	2709	));
			
  U2754	: Soma_AMA3_1 PORT MAP(
	A=> C(	2818	),
	B=>E(	2648	),
	Cin=> Carry( 	2753	),
	Cout=> Carry( 	2754	),
	S=> E(	2710	));
			
  U2755	: Soma_AMA3_1 PORT MAP(
	A=> C(	2819	),
	B=>E(	2649	),
	Cin=> Carry( 	2754	),
	Cout=> Carry( 	2755	),
	S=> E(	2711	));
			
  U2756	: Soma_AMA3_1 PORT MAP(
	A=> C(	2820	),
	B=>E(	2650	),
	Cin=> Carry( 	2755	),
	Cout=> Carry( 	2756	),
	S=> E(	2712	));
			
  U2757	: Soma_AMA3_1 PORT MAP(
	A=> C(	2821	),
	B=>E(	2651	),
	Cin=> Carry( 	2756	),
	Cout=> Carry( 	2757	),
	S=> E(	2713	));
			
  U2758	: Soma_AMA3_1 PORT MAP(
	A=> C(	2822	),
	B=>E(	2652	),
	Cin=> Carry( 	2757	),
	Cout=> Carry( 	2758	),
	S=> E(	2714	));
			
  U2759	: Soma_AMA3_1 PORT MAP(
	A=> C(	2823	),
	B=>E(	2653	),
	Cin=> Carry( 	2758	),
	Cout=> Carry( 	2759	),
	S=> E(	2715	));
			
  U2760	: Soma_AMA3_1 PORT MAP(
	A=> C(	2824	),
	B=>E(	2654	),
	Cin=> Carry( 	2759	),
	Cout=> Carry( 	2760	),
	S=> E(	2716	));
			
  U2761	: Soma_AMA3_1 PORT MAP(
	A=> C(	2825	),
	B=>E(	2655	),
	Cin=> Carry( 	2760	),
	Cout=> Carry( 	2761	),
	S=> E(	2717	));
			
  U2762	: Soma_AMA3_1 PORT MAP(
	A=> C(	2826	),
	B=>E(	2656	),
	Cin=> Carry( 	2761	),
	Cout=> Carry( 	2762	),
	S=> E(	2718	));
			
  U2763	: Soma_AMA3_1 PORT MAP(
	A=> C(	2827	),
	B=>E(	2657	),
	Cin=> Carry( 	2762	),
	Cout=> Carry( 	2763	),
	S=> E(	2719	));
			
  U2764	: Soma_AMA3_1 PORT MAP(
	A=> C(	2828	),
	B=>E(	2658	),
	Cin=> Carry( 	2763	),
	Cout=> Carry( 	2764	),
	S=> E(	2720	));
			
  U2765	: Soma_AMA3_1 PORT MAP(
	A=> C(	2829	),
	B=>E(	2659	),
	Cin=> Carry( 	2764	),
	Cout=> Carry( 	2765	),
	S=> E(	2721	));
			
  U2766	: Soma_AMA3_1 PORT MAP(
	A=> C(	2830	),
	B=>E(	2660	),
	Cin=> Carry( 	2765	),
	Cout=> Carry( 	2766	),
	S=> E(	2722	));
			
  U2767	: Soma_AMA3_1 PORT MAP(
	A=> C(	2831	),
	B=>E(	2661	),
	Cin=> Carry( 	2766	),
	Cout=> Carry( 	2767	),
	S=> E(	2723	));
			
  U2768	: Soma_AMA3_1 PORT MAP(
	A=> C(	2832	),
	B=>E(	2662	),
	Cin=> Carry( 	2767	),
	Cout=> Carry( 	2768	),
	S=> E(	2724	));
			
  U2769	: Soma_AMA3_1 PORT MAP(
	A=> C(	2833	),
	B=>E(	2663	),
	Cin=> Carry( 	2768	),
	Cout=> Carry( 	2769	),
	S=> E(	2725	));
			
  U2770	: Soma_AMA3_1 PORT MAP(
	A=> C(	2834	),
	B=>E(	2664	),
	Cin=> Carry( 	2769	),
	Cout=> Carry( 	2770	),
	S=> E(	2726	));
			
  U2771	: Soma_AMA3_1 PORT MAP(
	A=> C(	2835	),
	B=>E(	2665	),
	Cin=> Carry( 	2770	),
	Cout=> Carry( 	2771	),
	S=> E(	2727	));
			
  U2772	: Soma_AMA3_1 PORT MAP(
	A=> C(	2836	),
	B=>E(	2666	),
	Cin=> Carry( 	2771	),
	Cout=> Carry( 	2772	),
	S=> E(	2728	));
			
  U2773	: Soma_AMA3_1 PORT MAP(
	A=> C(	2837	),
	B=>E(	2667	),
	Cin=> Carry( 	2772	),
	Cout=> Carry( 	2773	),
	S=> E(	2729	));
			
  U2774	: Soma_AMA3_1 PORT MAP(
	A=> C(	2838	),
	B=>E(	2668	),
	Cin=> Carry( 	2773	),
	Cout=> Carry( 	2774	),
	S=> E(	2730	));
			
  U2775	: Soma_AMA3_1 PORT MAP(
	A=> C(	2839	),
	B=>E(	2669	),
	Cin=> Carry( 	2774	),
	Cout=> Carry( 	2775	),
	S=> E(	2731	));
			
  U2776	: Soma_AMA3_1 PORT MAP(
	A=> C(	2840	),
	B=>E(	2670	),
	Cin=> Carry( 	2775	),
	Cout=> Carry( 	2776	),
	S=> E(	2732	));
			
  U2777	: Soma_AMA3_1 PORT MAP(
	A=> C(	2841	),
	B=>E(	2671	),
	Cin=> Carry( 	2776	),
	Cout=> Carry( 	2777	),
	S=> E(	2733	));
			
  U2778	: Soma_AMA3_1 PORT MAP(
	A=> C(	2842	),
	B=>E(	2672	),
	Cin=> Carry( 	2777	),
	Cout=> Carry( 	2778	),
	S=> E(	2734	));
			
  U2779	: Soma_AMA3_1 PORT MAP(
	A=> C(	2843	),
	B=>E(	2673	),
	Cin=> Carry( 	2778	),
	Cout=> Carry( 	2779	),
	S=> E(	2735	));
			
  U2780	: Soma_AMA3_1 PORT MAP(
	A=> C(	2844	),
	B=>E(	2674	),
	Cin=> Carry( 	2779	),
	Cout=> Carry( 	2780	),
	S=> E(	2736	));
			
  U2781	: Soma_AMA3_1 PORT MAP(
	A=> C(	2845	),
	B=>E(	2675	),
	Cin=> Carry( 	2780	),
	Cout=> Carry( 	2781	),
	S=> E(	2737	));
			
  U2782	: Soma_AMA3_1 PORT MAP(
	A=> C(	2846	),
	B=>E(	2676	),
	Cin=> Carry( 	2781	),
	Cout=> Carry( 	2782	),
	S=> E(	2738	));
			
  U2783	: Soma_AMA3_1 PORT MAP(
	A=> C(	2847	),
	B=>E(	2677	),
	Cin=> Carry( 	2782	),
	Cout=> Carry( 	2783	),
	S=> E(	2739	));
			
  U2784	: Soma_AMA3_1 PORT MAP(
	A=> C(	2848	),
	B=>E(	2678	),
	Cin=> Carry( 	2783	),
	Cout=> Carry( 	2784	),
	S=> E(	2740	));
			
  U2785	: Soma_AMA3_1 PORT MAP(
	A=> C(	2849	),
	B=>E(	2679	),
	Cin=> Carry( 	2784	),
	Cout=> Carry( 	2785	),
	S=> E(	2741	));
			
  U2786	: Soma_AMA3_1 PORT MAP(
	A=> C(	2850	),
	B=>E(	2680	),
	Cin=> Carry( 	2785	),
	Cout=> Carry( 	2786	),
	S=> E(	2742	));
			
  U2787	: Soma_AMA3_1 PORT MAP(
	A=> C(	2851	),
	B=>E(	2681	),
	Cin=> Carry( 	2786	),
	Cout=> Carry( 	2787	),
	S=> E(	2743	));
			
  U2788	: Soma_AMA3_1 PORT MAP(
	A=> C(	2852	),
	B=>E(	2682	),
	Cin=> Carry( 	2787	),
	Cout=> Carry( 	2788	),
	S=> E(	2744	));
			
  U2789	: Soma_AMA3_1 PORT MAP(
	A=> C(	2853	),
	B=>E(	2683	),
	Cin=> Carry( 	2788	),
	Cout=> Carry( 	2789	),
	S=> E(	2745	));
			
  U2790	: Soma_AMA3_1 PORT MAP(
	A=> C(	2854	),
	B=>E(	2684	),
	Cin=> Carry( 	2789	),
	Cout=> Carry( 	2790	),
	S=> E(	2746	));
			
  U2791	: Soma_AMA3_1 PORT MAP(
	A=> C(	2855	),
	B=>E(	2685	),
	Cin=> Carry( 	2790	),
	Cout=> Carry( 	2791	),
	S=> E(	2747	));
			
  U2792	: Soma_AMA3_1 PORT MAP(
	A=> C(	2856	),
	B=>E(	2686	),
	Cin=> Carry( 	2791	),
	Cout=> Carry( 	2792	),
	S=> E(	2748	));
			
  U2793	: Soma_AMA3_1 PORT MAP(
	A=> C(	2857	),
	B=>E(	2687	),
	Cin=> Carry( 	2792	),
	Cout=> Carry( 	2793	),
	S=> E(	2749	));
			
  U2794	: Soma_AMA3_1 PORT MAP(
	A=> C(	2858	),
	B=>E(	2688	),
	Cin=> Carry( 	2793	),
	Cout=> Carry( 	2794	),
	S=> E(	2750	));
			
  U2795	: Soma_AMA3_1 PORT MAP(
	A=> C(	2859	),
	B=>E(	2689	),
	Cin=> Carry( 	2794	),
	Cout=> Carry( 	2795	),
	S=> E(	2751	));
			
  U2796	: Soma_AMA3_1 PORT MAP(
	A=> C(	2860	),
	B=>E(	2690	),
	Cin=> Carry( 	2795	),
	Cout=> Carry( 	2796	),
	S=> E(	2752	));
			
  U2797	: Soma_AMA3_1 PORT MAP(
	A=> C(	2861	),
	B=>E(	2691	),
	Cin=> Carry( 	2796	),
	Cout=> Carry( 	2797	),
	S=> E(	2753	));
			
  U2798	: Soma_AMA3_1 PORT MAP(
	A=> C(	2862	),
	B=>E(	2692	),
	Cin=> Carry( 	2797	),
	Cout=> Carry( 	2798	),
	S=> E(	2754	));
			
  U2799	: Soma_AMA3_1 PORT MAP(
	A=> C(	2863	),
	B=>E(	2693	),
	Cin=> Carry( 	2798	),
	Cout=> Carry( 	2799	),
	S=> E(	2755	));
			
  U2800	: Soma_AMA3_1 PORT MAP(
	A=> C(	2864	),
	B=>E(	2694	),
	Cin=> Carry( 	2799	),
	Cout=> Carry( 	2800	),
	S=> E(	2756	));
			
  U2801	: Soma_AMA3_1 PORT MAP(
	A=> C(	2865	),
	B=>E(	2695	),
	Cin=> Carry( 	2800	),
	Cout=> Carry( 	2801	),
	S=> E(	2757	));
			
  U2802	: Soma_AMA3_1 PORT MAP(
	A=> C(	2866	),
	B=>E(	2696	),
	Cin=> Carry( 	2801	),
	Cout=> Carry( 	2802	),
	S=> E(	2758	));
			
  U2803	: Soma_AMA3_1 PORT MAP(
	A=> C(	2867	),
	B=>E(	2697	),
	Cin=> Carry( 	2802	),
	Cout=> Carry( 	2803	),
	S=> E(	2759	));
			
  U2804	: Soma_AMA3_1 PORT MAP(
	A=> C(	2868	),
	B=>E(	2698	),
	Cin=> Carry( 	2803	),
	Cout=> Carry( 	2804	),
	S=> E(	2760	));
			
  U2805	: Soma_AMA3_1 PORT MAP(
	A=> C(	2869	),
	B=>E(	2699	),
	Cin=> Carry( 	2804	),
	Cout=> Carry( 	2805	),
	S=> E(	2761	));
			
  U2806	: Soma_AMA3_1 PORT MAP(
	A=> C(	2870	),
	B=>E(	2700	),
	Cin=> Carry( 	2805	),
	Cout=> Carry( 	2806	),
	S=> E(	2762	));
			
  U2807	: Soma_AMA3_1 PORT MAP(
	A=> C(	2871	),
	B=>E(	2701	),
	Cin=> Carry( 	2806	),
	Cout=> Carry( 	2807	),
	S=> E(	2763	));
			
  U2808	: Soma_AMA3_1 PORT MAP(
	A=> C(	2872	),
	B=>E(	2702	),
	Cin=> Carry( 	2807	),
	Cout=> Carry( 	2808	),
	S=> E(	2764	));
			
  U2809	: Soma_AMA3_1 PORT MAP(
	A=> C(	2873	),
	B=>E(	2703	),
	Cin=> Carry( 	2808	),
	Cout=> Carry( 	2809	),
	S=> E(	2765	));
			
  U2810	: Soma_AMA3_1 PORT MAP(
	A=> C(	2874	),
	B=>E(	2704	),
	Cin=> Carry( 	2809	),
	Cout=> Carry( 	2810	),
	S=> E(	2766	));
			
  U2811	: Soma_AMA3_1 PORT MAP(
	A=> C(	2875	),
	B=>E(	2705	),
	Cin=> Carry( 	2810	),
	Cout=> Carry( 	2811	),
	S=> E(	2767	));
			
  U2812	: Soma_AMA3_1 PORT MAP(
	A=> C(	2876	),
	B=>E(	2706	),
	Cin=> Carry( 	2811	),
	Cout=> Carry( 	2812	),
	S=> E(	2768	));
			
  U2813	: Soma_AMA3_1 PORT MAP(
	A=> C(	2877	),
	B=>E(	2707	),
	Cin=> Carry( 	2812	),
	Cout=> Carry( 	2813	),
	S=> E(	2769	));
			
  U2814	: Soma_AMA3_1 PORT MAP(
	A=> C(	2878	),
	B=>E(	2708	),
	Cin=> Carry( 	2813	),
	Cout=> Carry( 	2814	),
	S=> E(	2770	));
			
  U2815	: Soma_AMA3_1 PORT MAP(
	A=> C(	2879	),
	B=>Carry(	2751	),
	Cin=> Carry( 	2814	),
	Cout=> Carry( 	2815	),
	S=> E(	2771	));


			
  U2816	: Soma_AMA3_1 PORT MAP(
	A=> C(	2880	),
	B=>E(	2709	),
	Cin=> '0'	,
	Cout=> Carry( 	2816	),
	S=> R(	45	));
			
  U2817	: Soma_AMA3_1 PORT MAP(
	A=> C(	2881	),
	B=>E(	2710	),
	Cin=> Carry( 	2816	),
	Cout=> Carry( 	2817	),
	S=> E(	2772	));
			
  U2818	: Soma_AMA3_1 PORT MAP(
	A=> C(	2882	),
	B=>E(	2711	),
	Cin=> Carry( 	2817	),
	Cout=> Carry( 	2818	),
	S=> E(	2773	));
			
  U2819	: Soma_AMA3_1 PORT MAP(
	A=> C(	2883	),
	B=>E(	2712	),
	Cin=> Carry( 	2818	),
	Cout=> Carry( 	2819	),
	S=> E(	2774	));
			
  U2820	: Soma_AMA3_1 PORT MAP(
	A=> C(	2884	),
	B=>E(	2713	),
	Cin=> Carry( 	2819	),
	Cout=> Carry( 	2820	),
	S=> E(	2775	));
			
  U2821	: Soma_AMA3_1 PORT MAP(
	A=> C(	2885	),
	B=>E(	2714	),
	Cin=> Carry( 	2820	),
	Cout=> Carry( 	2821	),
	S=> E(	2776	));
			
  U2822	: Soma_AMA3_1 PORT MAP(
	A=> C(	2886	),
	B=>E(	2715	),
	Cin=> Carry( 	2821	),
	Cout=> Carry( 	2822	),
	S=> E(	2777	));
			
  U2823	: Soma_AMA3_1 PORT MAP(
	A=> C(	2887	),
	B=>E(	2716	),
	Cin=> Carry( 	2822	),
	Cout=> Carry( 	2823	),
	S=> E(	2778	));
			
  U2824	: Soma_AMA3_1 PORT MAP(
	A=> C(	2888	),
	B=>E(	2717	),
	Cin=> Carry( 	2823	),
	Cout=> Carry( 	2824	),
	S=> E(	2779	));
			
  U2825	: Soma_AMA3_1 PORT MAP(
	A=> C(	2889	),
	B=>E(	2718	),
	Cin=> Carry( 	2824	),
	Cout=> Carry( 	2825	),
	S=> E(	2780	));
			
  U2826	: Soma_AMA3_1 PORT MAP(
	A=> C(	2890	),
	B=>E(	2719	),
	Cin=> Carry( 	2825	),
	Cout=> Carry( 	2826	),
	S=> E(	2781	));
			
  U2827	: Soma_AMA3_1 PORT MAP(
	A=> C(	2891	),
	B=>E(	2720	),
	Cin=> Carry( 	2826	),
	Cout=> Carry( 	2827	),
	S=> E(	2782	));
			
  U2828	: Soma_AMA3_1 PORT MAP(
	A=> C(	2892	),
	B=>E(	2721	),
	Cin=> Carry( 	2827	),
	Cout=> Carry( 	2828	),
	S=> E(	2783	));
			
  U2829	: Soma_AMA3_1 PORT MAP(
	A=> C(	2893	),
	B=>E(	2722	),
	Cin=> Carry( 	2828	),
	Cout=> Carry( 	2829	),
	S=> E(	2784	));
			
  U2830	: Soma_AMA3_1 PORT MAP(
	A=> C(	2894	),
	B=>E(	2723	),
	Cin=> Carry( 	2829	),
	Cout=> Carry( 	2830	),
	S=> E(	2785	));
			
  U2831	: Soma_AMA3_1 PORT MAP(
	A=> C(	2895	),
	B=>E(	2724	),
	Cin=> Carry( 	2830	),
	Cout=> Carry( 	2831	),
	S=> E(	2786	));
			
  U2832	: Soma_AMA3_1 PORT MAP(
	A=> C(	2896	),
	B=>E(	2725	),
	Cin=> Carry( 	2831	),
	Cout=> Carry( 	2832	),
	S=> E(	2787	));
			
  U2833	: Soma_AMA3_1 PORT MAP(
	A=> C(	2897	),
	B=>E(	2726	),
	Cin=> Carry( 	2832	),
	Cout=> Carry( 	2833	),
	S=> E(	2788	));
			
  U2834	: Soma_AMA3_1 PORT MAP(
	A=> C(	2898	),
	B=>E(	2727	),
	Cin=> Carry( 	2833	),
	Cout=> Carry( 	2834	),
	S=> E(	2789	));
			
  U2835	: Soma_AMA3_1 PORT MAP(
	A=> C(	2899	),
	B=>E(	2728	),
	Cin=> Carry( 	2834	),
	Cout=> Carry( 	2835	),
	S=> E(	2790	));
			
  U2836	: Soma_AMA3_1 PORT MAP(
	A=> C(	2900	),
	B=>E(	2729	),
	Cin=> Carry( 	2835	),
	Cout=> Carry( 	2836	),
	S=> E(	2791	));
			
  U2837	: Soma_AMA3_1 PORT MAP(
	A=> C(	2901	),
	B=>E(	2730	),
	Cin=> Carry( 	2836	),
	Cout=> Carry( 	2837	),
	S=> E(	2792	));
			
  U2838	: Soma_AMA3_1 PORT MAP(
	A=> C(	2902	),
	B=>E(	2731	),
	Cin=> Carry( 	2837	),
	Cout=> Carry( 	2838	),
	S=> E(	2793	));
			
  U2839	: Soma_AMA3_1 PORT MAP(
	A=> C(	2903	),
	B=>E(	2732	),
	Cin=> Carry( 	2838	),
	Cout=> Carry( 	2839	),
	S=> E(	2794	));
			
  U2840	: Soma_AMA3_1 PORT MAP(
	A=> C(	2904	),
	B=>E(	2733	),
	Cin=> Carry( 	2839	),
	Cout=> Carry( 	2840	),
	S=> E(	2795	));
			
  U2841	: Soma_AMA3_1 PORT MAP(
	A=> C(	2905	),
	B=>E(	2734	),
	Cin=> Carry( 	2840	),
	Cout=> Carry( 	2841	),
	S=> E(	2796	));
			
  U2842	: Soma_AMA3_1 PORT MAP(
	A=> C(	2906	),
	B=>E(	2735	),
	Cin=> Carry( 	2841	),
	Cout=> Carry( 	2842	),
	S=> E(	2797	));
			
  U2843	: Soma_AMA3_1 PORT MAP(
	A=> C(	2907	),
	B=>E(	2736	),
	Cin=> Carry( 	2842	),
	Cout=> Carry( 	2843	),
	S=> E(	2798	));
			
  U2844	: Soma_AMA3_1 PORT MAP(
	A=> C(	2908	),
	B=>E(	2737	),
	Cin=> Carry( 	2843	),
	Cout=> Carry( 	2844	),
	S=> E(	2799	));
			
  U2845	: Soma_AMA3_1 PORT MAP(
	A=> C(	2909	),
	B=>E(	2738	),
	Cin=> Carry( 	2844	),
	Cout=> Carry( 	2845	),
	S=> E(	2800	));
			
  U2846	: Soma_AMA3_1 PORT MAP(
	A=> C(	2910	),
	B=>E(	2739	),
	Cin=> Carry( 	2845	),
	Cout=> Carry( 	2846	),
	S=> E(	2801	));
			
  U2847	: Soma_AMA3_1 PORT MAP(
	A=> C(	2911	),
	B=>E(	2740	),
	Cin=> Carry( 	2846	),
	Cout=> Carry( 	2847	),
	S=> E(	2802	));
			
  U2848	: Soma_AMA3_1 PORT MAP(
	A=> C(	2912	),
	B=>E(	2741	),
	Cin=> Carry( 	2847	),
	Cout=> Carry( 	2848	),
	S=> E(	2803	));
			
  U2849	: Soma_AMA3_1 PORT MAP(
	A=> C(	2913	),
	B=>E(	2742	),
	Cin=> Carry( 	2848	),
	Cout=> Carry( 	2849	),
	S=> E(	2804	));
			
  U2850	: Soma_AMA3_1 PORT MAP(
	A=> C(	2914	),
	B=>E(	2743	),
	Cin=> Carry( 	2849	),
	Cout=> Carry( 	2850	),
	S=> E(	2805	));
			
  U2851	: Soma_AMA3_1 PORT MAP(
	A=> C(	2915	),
	B=>E(	2744	),
	Cin=> Carry( 	2850	),
	Cout=> Carry( 	2851	),
	S=> E(	2806	));
			
  U2852	: Soma_AMA3_1 PORT MAP(
	A=> C(	2916	),
	B=>E(	2745	),
	Cin=> Carry( 	2851	),
	Cout=> Carry( 	2852	),
	S=> E(	2807	));
			
  U2853	: Soma_AMA3_1 PORT MAP(
	A=> C(	2917	),
	B=>E(	2746	),
	Cin=> Carry( 	2852	),
	Cout=> Carry( 	2853	),
	S=> E(	2808	));
			
  U2854	: Soma_AMA3_1 PORT MAP(
	A=> C(	2918	),
	B=>E(	2747	),
	Cin=> Carry( 	2853	),
	Cout=> Carry( 	2854	),
	S=> E(	2809	));
			
  U2855	: Soma_AMA3_1 PORT MAP(
	A=> C(	2919	),
	B=>E(	2748	),
	Cin=> Carry( 	2854	),
	Cout=> Carry( 	2855	),
	S=> E(	2810	));
			
  U2856	: Soma_AMA3_1 PORT MAP(
	A=> C(	2920	),
	B=>E(	2749	),
	Cin=> Carry( 	2855	),
	Cout=> Carry( 	2856	),
	S=> E(	2811	));
			
  U2857	: Soma_AMA3_1 PORT MAP(
	A=> C(	2921	),
	B=>E(	2750	),
	Cin=> Carry( 	2856	),
	Cout=> Carry( 	2857	),
	S=> E(	2812	));
			
  U2858	: Soma_AMA3_1 PORT MAP(
	A=> C(	2922	),
	B=>E(	2751	),
	Cin=> Carry( 	2857	),
	Cout=> Carry( 	2858	),
	S=> E(	2813	));
			
  U2859	: Soma_AMA3_1 PORT MAP(
	A=> C(	2923	),
	B=>E(	2752	),
	Cin=> Carry( 	2858	),
	Cout=> Carry( 	2859	),
	S=> E(	2814	));
			
  U2860	: Soma_AMA3_1 PORT MAP(
	A=> C(	2924	),
	B=>E(	2753	),
	Cin=> Carry( 	2859	),
	Cout=> Carry( 	2860	),
	S=> E(	2815	));
			
  U2861	: Soma_AMA3_1 PORT MAP(
	A=> C(	2925	),
	B=>E(	2754	),
	Cin=> Carry( 	2860	),
	Cout=> Carry( 	2861	),
	S=> E(	2816	));
			
  U2862	: Soma_AMA3_1 PORT MAP(
	A=> C(	2926	),
	B=>E(	2755	),
	Cin=> Carry( 	2861	),
	Cout=> Carry( 	2862	),
	S=> E(	2817	));
			
  U2863	: Soma_AMA3_1 PORT MAP(
	A=> C(	2927	),
	B=>E(	2756	),
	Cin=> Carry( 	2862	),
	Cout=> Carry( 	2863	),
	S=> E(	2818	));
			
  U2864	: Soma_AMA3_1 PORT MAP(
	A=> C(	2928	),
	B=>E(	2757	),
	Cin=> Carry( 	2863	),
	Cout=> Carry( 	2864	),
	S=> E(	2819	));
			
  U2865	: Soma_AMA3_1 PORT MAP(
	A=> C(	2929	),
	B=>E(	2758	),
	Cin=> Carry( 	2864	),
	Cout=> Carry( 	2865	),
	S=> E(	2820	));
			
  U2866	: Soma_AMA3_1 PORT MAP(
	A=> C(	2930	),
	B=>E(	2759	),
	Cin=> Carry( 	2865	),
	Cout=> Carry( 	2866	),
	S=> E(	2821	));
			
  U2867	: Soma_AMA3_1 PORT MAP(
	A=> C(	2931	),
	B=>E(	2760	),
	Cin=> Carry( 	2866	),
	Cout=> Carry( 	2867	),
	S=> E(	2822	));
			
  U2868	: Soma_AMA3_1 PORT MAP(
	A=> C(	2932	),
	B=>E(	2761	),
	Cin=> Carry( 	2867	),
	Cout=> Carry( 	2868	),
	S=> E(	2823	));
			
  U2869	: Soma_AMA3_1 PORT MAP(
	A=> C(	2933	),
	B=>E(	2762	),
	Cin=> Carry( 	2868	),
	Cout=> Carry( 	2869	),
	S=> E(	2824	));
			
  U2870	: Soma_AMA3_1 PORT MAP(
	A=> C(	2934	),
	B=>E(	2763	),
	Cin=> Carry( 	2869	),
	Cout=> Carry( 	2870	),
	S=> E(	2825	));
			
  U2871	: Soma_AMA3_1 PORT MAP(
	A=> C(	2935	),
	B=>E(	2764	),
	Cin=> Carry( 	2870	),
	Cout=> Carry( 	2871	),
	S=> E(	2826	));
			
  U2872	: Soma_AMA3_1 PORT MAP(
	A=> C(	2936	),
	B=>E(	2765	),
	Cin=> Carry( 	2871	),
	Cout=> Carry( 	2872	),
	S=> E(	2827	));
			
  U2873	: Soma_AMA3_1 PORT MAP(
	A=> C(	2937	),
	B=>E(	2766	),
	Cin=> Carry( 	2872	),
	Cout=> Carry( 	2873	),
	S=> E(	2828	));
			
  U2874	: Soma_AMA3_1 PORT MAP(
	A=> C(	2938	),
	B=>E(	2767	),
	Cin=> Carry( 	2873	),
	Cout=> Carry( 	2874	),
	S=> E(	2829	));
			
  U2875	: Soma_AMA3_1 PORT MAP(
	A=> C(	2939	),
	B=>E(	2768	),
	Cin=> Carry( 	2874	),
	Cout=> Carry( 	2875	),
	S=> E(	2830	));
			
  U2876	: Soma_AMA3_1 PORT MAP(
	A=> C(	2940	),
	B=>E(	2769	),
	Cin=> Carry( 	2875	),
	Cout=> Carry( 	2876	),
	S=> E(	2831	));
			
  U2877	: Soma_AMA3_1 PORT MAP(
	A=> C(	2941	),
	B=>E(	2770	),
	Cin=> Carry( 	2876	),
	Cout=> Carry( 	2877	),
	S=> E(	2832	));
			
  U2878	: Soma_AMA3_1 PORT MAP(
	A=> C(	2942	),
	B=>E(	2771	),
	Cin=> Carry( 	2877	),
	Cout=> Carry( 	2878	),
	S=> E(	2833	));
			
  U2879	: Soma_AMA3_1 PORT MAP(
	A=> C(	2943	),
	B=>Carry(	2815	),
	Cin=> Carry( 	2878	),
	Cout=> Carry( 	2879	),
	S=> E(	2834	));

			
  U2880	: Soma_AMA3_1 PORT MAP(
	A=> C(	2944	),
	B=>E(	2772	),
	Cin=> '0'	,
	Cout=> Carry( 	2880	),
	S=> R(	46	));
			
  U2881	: Soma_AMA3_1 PORT MAP(
	A=> C(	2945	),
	B=>E(	2773	),
	Cin=> Carry( 	2880	),
	Cout=> Carry( 	2881	),
	S=> E(	2835	));
			
  U2882	: Soma_AMA3_1 PORT MAP(
	A=> C(	2946	),
	B=>E(	2774	),
	Cin=> Carry( 	2881	),
	Cout=> Carry( 	2882	),
	S=> E(	2836	));
			
  U2883	: Soma_AMA3_1 PORT MAP(
	A=> C(	2947	),
	B=>E(	2775	),
	Cin=> Carry( 	2882	),
	Cout=> Carry( 	2883	),
	S=> E(	2837	));
			
  U2884	: Soma_AMA3_1 PORT MAP(
	A=> C(	2948	),
	B=>E(	2776	),
	Cin=> Carry( 	2883	),
	Cout=> Carry( 	2884	),
	S=> E(	2838	));
			
  U2885	: Soma_AMA3_1 PORT MAP(
	A=> C(	2949	),
	B=>E(	2777	),
	Cin=> Carry( 	2884	),
	Cout=> Carry( 	2885	),
	S=> E(	2839	));
			
  U2886	: Soma_AMA3_1 PORT MAP(
	A=> C(	2950	),
	B=>E(	2778	),
	Cin=> Carry( 	2885	),
	Cout=> Carry( 	2886	),
	S=> E(	2840	));
			
  U2887	: Soma_AMA3_1 PORT MAP(
	A=> C(	2951	),
	B=>E(	2779	),
	Cin=> Carry( 	2886	),
	Cout=> Carry( 	2887	),
	S=> E(	2841	));
			
  U2888	: Soma_AMA3_1 PORT MAP(
	A=> C(	2952	),
	B=>E(	2780	),
	Cin=> Carry( 	2887	),
	Cout=> Carry( 	2888	),
	S=> E(	2842	));
			
  U2889	: Soma_AMA3_1 PORT MAP(
	A=> C(	2953	),
	B=>E(	2781	),
	Cin=> Carry( 	2888	),
	Cout=> Carry( 	2889	),
	S=> E(	2843	));
			
  U2890	: Soma_AMA3_1 PORT MAP(
	A=> C(	2954	),
	B=>E(	2782	),
	Cin=> Carry( 	2889	),
	Cout=> Carry( 	2890	),
	S=> E(	2844	));
			
  U2891	: Soma_AMA3_1 PORT MAP(
	A=> C(	2955	),
	B=>E(	2783	),
	Cin=> Carry( 	2890	),
	Cout=> Carry( 	2891	),
	S=> E(	2845	));
			
  U2892	: Soma_AMA3_1 PORT MAP(
	A=> C(	2956	),
	B=>E(	2784	),
	Cin=> Carry( 	2891	),
	Cout=> Carry( 	2892	),
	S=> E(	2846	));
			
  U2893	: Soma_AMA3_1 PORT MAP(
	A=> C(	2957	),
	B=>E(	2785	),
	Cin=> Carry( 	2892	),
	Cout=> Carry( 	2893	),
	S=> E(	2847	));
			
  U2894	: Soma_AMA3_1 PORT MAP(
	A=> C(	2958	),
	B=>E(	2786	),
	Cin=> Carry( 	2893	),
	Cout=> Carry( 	2894	),
	S=> E(	2848	));
			
  U2895	: Soma_AMA3_1 PORT MAP(
	A=> C(	2959	),
	B=>E(	2787	),
	Cin=> Carry( 	2894	),
	Cout=> Carry( 	2895	),
	S=> E(	2849	));
			
  U2896	: Soma_AMA3_1 PORT MAP(
	A=> C(	2960	),
	B=>E(	2788	),
	Cin=> Carry( 	2895	),
	Cout=> Carry( 	2896	),
	S=> E(	2850	));
			
  U2897	: Soma_AMA3_1 PORT MAP(
	A=> C(	2961	),
	B=>E(	2789	),
	Cin=> Carry( 	2896	),
	Cout=> Carry( 	2897	),
	S=> E(	2851	));
			
  U2898	: Soma_AMA3_1 PORT MAP(
	A=> C(	2962	),
	B=>E(	2790	),
	Cin=> Carry( 	2897	),
	Cout=> Carry( 	2898	),
	S=> E(	2852	));
			
  U2899	: Soma_AMA3_1 PORT MAP(
	A=> C(	2963	),
	B=>E(	2791	),
	Cin=> Carry( 	2898	),
	Cout=> Carry( 	2899	),
	S=> E(	2853	));
			
  U2900	: Soma_AMA3_1 PORT MAP(
	A=> C(	2964	),
	B=>E(	2792	),
	Cin=> Carry( 	2899	),
	Cout=> Carry( 	2900	),
	S=> E(	2854	));
			
  U2901	: Soma_AMA3_1 PORT MAP(
	A=> C(	2965	),
	B=>E(	2793	),
	Cin=> Carry( 	2900	),
	Cout=> Carry( 	2901	),
	S=> E(	2855	));
			
  U2902	: Soma_AMA3_1 PORT MAP(
	A=> C(	2966	),
	B=>E(	2794	),
	Cin=> Carry( 	2901	),
	Cout=> Carry( 	2902	),
	S=> E(	2856	));
			
  U2903	: Soma_AMA3_1 PORT MAP(
	A=> C(	2967	),
	B=>E(	2795	),
	Cin=> Carry( 	2902	),
	Cout=> Carry( 	2903	),
	S=> E(	2857	));
			
  U2904	: Soma_AMA3_1 PORT MAP(
	A=> C(	2968	),
	B=>E(	2796	),
	Cin=> Carry( 	2903	),
	Cout=> Carry( 	2904	),
	S=> E(	2858	));
			
  U2905	: Soma_AMA3_1 PORT MAP(
	A=> C(	2969	),
	B=>E(	2797	),
	Cin=> Carry( 	2904	),
	Cout=> Carry( 	2905	),
	S=> E(	2859	));
			
  U2906	: Soma_AMA3_1 PORT MAP(
	A=> C(	2970	),
	B=>E(	2798	),
	Cin=> Carry( 	2905	),
	Cout=> Carry( 	2906	),
	S=> E(	2860	));
			
  U2907	: Soma_AMA3_1 PORT MAP(
	A=> C(	2971	),
	B=>E(	2799	),
	Cin=> Carry( 	2906	),
	Cout=> Carry( 	2907	),
	S=> E(	2861	));
			
  U2908	: Soma_AMA3_1 PORT MAP(
	A=> C(	2972	),
	B=>E(	2800	),
	Cin=> Carry( 	2907	),
	Cout=> Carry( 	2908	),
	S=> E(	2862	));
			
  U2909	: Soma_AMA3_1 PORT MAP(
	A=> C(	2973	),
	B=>E(	2801	),
	Cin=> Carry( 	2908	),
	Cout=> Carry( 	2909	),
	S=> E(	2863	));
			
  U2910	: Soma_AMA3_1 PORT MAP(
	A=> C(	2974	),
	B=>E(	2802	),
	Cin=> Carry( 	2909	),
	Cout=> Carry( 	2910	),
	S=> E(	2864	));
			
  U2911	: Soma_AMA3_1 PORT MAP(
	A=> C(	2975	),
	B=>E(	2803	),
	Cin=> Carry( 	2910	),
	Cout=> Carry( 	2911	),
	S=> E(	2865	));
			
  U2912	: Soma_AMA3_1 PORT MAP(
	A=> C(	2976	),
	B=>E(	2804	),
	Cin=> Carry( 	2911	),
	Cout=> Carry( 	2912	),
	S=> E(	2866	));
			
  U2913	: Soma_AMA3_1 PORT MAP(
	A=> C(	2977	),
	B=>E(	2805	),
	Cin=> Carry( 	2912	),
	Cout=> Carry( 	2913	),
	S=> E(	2867	));
			
  U2914	: Soma_AMA3_1 PORT MAP(
	A=> C(	2978	),
	B=>E(	2806	),
	Cin=> Carry( 	2913	),
	Cout=> Carry( 	2914	),
	S=> E(	2868	));
			
  U2915	: Soma_AMA3_1 PORT MAP(
	A=> C(	2979	),
	B=>E(	2807	),
	Cin=> Carry( 	2914	),
	Cout=> Carry( 	2915	),
	S=> E(	2869	));
			
  U2916	: Soma_AMA3_1 PORT MAP(
	A=> C(	2980	),
	B=>E(	2808	),
	Cin=> Carry( 	2915	),
	Cout=> Carry( 	2916	),
	S=> E(	2870	));
			
  U2917	: Soma_AMA3_1 PORT MAP(
	A=> C(	2981	),
	B=>E(	2809	),
	Cin=> Carry( 	2916	),
	Cout=> Carry( 	2917	),
	S=> E(	2871	));
			
  U2918	: Soma_AMA3_1 PORT MAP(
	A=> C(	2982	),
	B=>E(	2810	),
	Cin=> Carry( 	2917	),
	Cout=> Carry( 	2918	),
	S=> E(	2872	));
			
  U2919	: Soma_AMA3_1 PORT MAP(
	A=> C(	2983	),
	B=>E(	2811	),
	Cin=> Carry( 	2918	),
	Cout=> Carry( 	2919	),
	S=> E(	2873	));
			
  U2920	: Soma_AMA3_1 PORT MAP(
	A=> C(	2984	),
	B=>E(	2812	),
	Cin=> Carry( 	2919	),
	Cout=> Carry( 	2920	),
	S=> E(	2874	));
			
  U2921	: Soma_AMA3_1 PORT MAP(
	A=> C(	2985	),
	B=>E(	2813	),
	Cin=> Carry( 	2920	),
	Cout=> Carry( 	2921	),
	S=> E(	2875	));
			
  U2922	: Soma_AMA3_1 PORT MAP(
	A=> C(	2986	),
	B=>E(	2814	),
	Cin=> Carry( 	2921	),
	Cout=> Carry( 	2922	),
	S=> E(	2876	));
			
  U2923	: Soma_AMA3_1 PORT MAP(
	A=> C(	2987	),
	B=>E(	2815	),
	Cin=> Carry( 	2922	),
	Cout=> Carry( 	2923	),
	S=> E(	2877	));
			
  U2924	: Soma_AMA3_1 PORT MAP(
	A=> C(	2988	),
	B=>E(	2816	),
	Cin=> Carry( 	2923	),
	Cout=> Carry( 	2924	),
	S=> E(	2878	));
			
  U2925	: Soma_AMA3_1 PORT MAP(
	A=> C(	2989	),
	B=>E(	2817	),
	Cin=> Carry( 	2924	),
	Cout=> Carry( 	2925	),
	S=> E(	2879	));
			
  U2926	: Soma_AMA3_1 PORT MAP(
	A=> C(	2990	),
	B=>E(	2818	),
	Cin=> Carry( 	2925	),
	Cout=> Carry( 	2926	),
	S=> E(	2880	));
			
  U2927	: Soma_AMA3_1 PORT MAP(
	A=> C(	2991	),
	B=>E(	2819	),
	Cin=> Carry( 	2926	),
	Cout=> Carry( 	2927	),
	S=> E(	2881	));
			
  U2928	: Soma_AMA3_1 PORT MAP(
	A=> C(	2992	),
	B=>E(	2820	),
	Cin=> Carry( 	2927	),
	Cout=> Carry( 	2928	),
	S=> E(	2882	));
			
  U2929	: Soma_AMA3_1 PORT MAP(
	A=> C(	2993	),
	B=>E(	2821	),
	Cin=> Carry( 	2928	),
	Cout=> Carry( 	2929	),
	S=> E(	2883	));
			
  U2930	: Soma_AMA3_1 PORT MAP(
	A=> C(	2994	),
	B=>E(	2822	),
	Cin=> Carry( 	2929	),
	Cout=> Carry( 	2930	),
	S=> E(	2884	));
			
  U2931	: Soma_AMA3_1 PORT MAP(
	A=> C(	2995	),
	B=>E(	2823	),
	Cin=> Carry( 	2930	),
	Cout=> Carry( 	2931	),
	S=> E(	2885	));
			
  U2932	: Soma_AMA3_1 PORT MAP(
	A=> C(	2996	),
	B=>E(	2824	),
	Cin=> Carry( 	2931	),
	Cout=> Carry( 	2932	),
	S=> E(	2886	));
			
  U2933	: Soma_AMA3_1 PORT MAP(
	A=> C(	2997	),
	B=>E(	2825	),
	Cin=> Carry( 	2932	),
	Cout=> Carry( 	2933	),
	S=> E(	2887	));
			
  U2934	: Soma_AMA3_1 PORT MAP(
	A=> C(	2998	),
	B=>E(	2826	),
	Cin=> Carry( 	2933	),
	Cout=> Carry( 	2934	),
	S=> E(	2888	));
			
  U2935	: Soma_AMA3_1 PORT MAP(
	A=> C(	2999	),
	B=>E(	2827	),
	Cin=> Carry( 	2934	),
	Cout=> Carry( 	2935	),
	S=> E(	2889	));
			
  U2936	: Soma_AMA3_1 PORT MAP(
	A=> C(	3000	),
	B=>E(	2828	),
	Cin=> Carry( 	2935	),
	Cout=> Carry( 	2936	),
	S=> E(	2890	));
			
  U2937	: Soma_AMA3_1 PORT MAP(
	A=> C(	3001	),
	B=>E(	2829	),
	Cin=> Carry( 	2936	),
	Cout=> Carry( 	2937	),
	S=> E(	2891	));
			
  U2938	: Soma_AMA3_1 PORT MAP(
	A=> C(	3002	),
	B=>E(	2830	),
	Cin=> Carry( 	2937	),
	Cout=> Carry( 	2938	),
	S=> E(	2892	));
			
  U2939	: Soma_AMA3_1 PORT MAP(
	A=> C(	3003	),
	B=>E(	2831	),
	Cin=> Carry( 	2938	),
	Cout=> Carry( 	2939	),
	S=> E(	2893	));
			
  U2940	: Soma_AMA3_1 PORT MAP(
	A=> C(	3004	),
	B=>E(	2832	),
	Cin=> Carry( 	2939	),
	Cout=> Carry( 	2940	),
	S=> E(	2894	));
			
  U2941	: Soma_AMA3_1 PORT MAP(
	A=> C(	3005	),
	B=>E(	2833	),
	Cin=> Carry( 	2940	),
	Cout=> Carry( 	2941	),
	S=> E(	2895	));
			
  U2942	: Soma_AMA3_1 PORT MAP(
	A=> C(	3006	),
	B=>E(	2834	),
	Cin=> Carry( 	2941	),
	Cout=> Carry( 	2942	),
	S=> E(	2896	));
			
  U2943	: Soma_AMA3_1 PORT MAP(
	A=> C(	3007	),
	B=>Carry(	2879	),
	Cin=> Carry( 	2942	),
	Cout=> Carry( 	2943	),
	S=> E(	2897	));

			
  U2944	: Soma_AMA3_1 PORT MAP(
	A=> C(	3008	),
	B=>E(	2835	),
	Cin=> '0'	,
	Cout=> Carry( 	2944	),
	S=> R(	47	));
			
  U2945	: Soma_AMA3_1 PORT MAP(
	A=> C(	3009	),
	B=>E(	2836	),
	Cin=> Carry( 	2944	),
	Cout=> Carry( 	2945	),
	S=> E(	2898	));
			
  U2946	: Soma_AMA3_1 PORT MAP(
	A=> C(	3010	),
	B=>E(	2837	),
	Cin=> Carry( 	2945	),
	Cout=> Carry( 	2946	),
	S=> E(	2899	));
			
  U2947	: Soma_AMA3_1 PORT MAP(
	A=> C(	3011	),
	B=>E(	2838	),
	Cin=> Carry( 	2946	),
	Cout=> Carry( 	2947	),
	S=> E(	2900	));
			
  U2948	: Soma_AMA3_1 PORT MAP(
	A=> C(	3012	),
	B=>E(	2839	),
	Cin=> Carry( 	2947	),
	Cout=> Carry( 	2948	),
	S=> E(	2901	));
			
  U2949	: Soma_AMA3_1 PORT MAP(
	A=> C(	3013	),
	B=>E(	2840	),
	Cin=> Carry( 	2948	),
	Cout=> Carry( 	2949	),
	S=> E(	2902	));
			
  U2950	: Soma_AMA3_1 PORT MAP(
	A=> C(	3014	),
	B=>E(	2841	),
	Cin=> Carry( 	2949	),
	Cout=> Carry( 	2950	),
	S=> E(	2903	));
			
  U2951	: Soma_AMA3_1 PORT MAP(
	A=> C(	3015	),
	B=>E(	2842	),
	Cin=> Carry( 	2950	),
	Cout=> Carry( 	2951	),
	S=> E(	2904	));
			
  U2952	: Soma_AMA3_1 PORT MAP(
	A=> C(	3016	),
	B=>E(	2843	),
	Cin=> Carry( 	2951	),
	Cout=> Carry( 	2952	),
	S=> E(	2905	));
			
  U2953	: Soma_AMA3_1 PORT MAP(
	A=> C(	3017	),
	B=>E(	2844	),
	Cin=> Carry( 	2952	),
	Cout=> Carry( 	2953	),
	S=> E(	2906	));
			
  U2954	: Soma_AMA3_1 PORT MAP(
	A=> C(	3018	),
	B=>E(	2845	),
	Cin=> Carry( 	2953	),
	Cout=> Carry( 	2954	),
	S=> E(	2907	));
			
  U2955	: Soma_AMA3_1 PORT MAP(
	A=> C(	3019	),
	B=>E(	2846	),
	Cin=> Carry( 	2954	),
	Cout=> Carry( 	2955	),
	S=> E(	2908	));
			
  U2956	: Soma_AMA3_1 PORT MAP(
	A=> C(	3020	),
	B=>E(	2847	),
	Cin=> Carry( 	2955	),
	Cout=> Carry( 	2956	),
	S=> E(	2909	));
			
  U2957	: Soma_AMA3_1 PORT MAP(
	A=> C(	3021	),
	B=>E(	2848	),
	Cin=> Carry( 	2956	),
	Cout=> Carry( 	2957	),
	S=> E(	2910	));
			
  U2958	: Soma_AMA3_1 PORT MAP(
	A=> C(	3022	),
	B=>E(	2849	),
	Cin=> Carry( 	2957	),
	Cout=> Carry( 	2958	),
	S=> E(	2911	));
			
  U2959	: Soma_AMA3_1 PORT MAP(
	A=> C(	3023	),
	B=>E(	2850	),
	Cin=> Carry( 	2958	),
	Cout=> Carry( 	2959	),
	S=> E(	2912	));
			
  U2960	: Soma_AMA3_1 PORT MAP(
	A=> C(	3024	),
	B=>E(	2851	),
	Cin=> Carry( 	2959	),
	Cout=> Carry( 	2960	),
	S=> E(	2913	));
			
  U2961	: Soma_AMA3_1 PORT MAP(
	A=> C(	3025	),
	B=>E(	2852	),
	Cin=> Carry( 	2960	),
	Cout=> Carry( 	2961	),
	S=> E(	2914	));
			
  U2962	: Soma_AMA3_1 PORT MAP(
	A=> C(	3026	),
	B=>E(	2853	),
	Cin=> Carry( 	2961	),
	Cout=> Carry( 	2962	),
	S=> E(	2915	));
			
  U2963	: Soma_AMA3_1 PORT MAP(
	A=> C(	3027	),
	B=>E(	2854	),
	Cin=> Carry( 	2962	),
	Cout=> Carry( 	2963	),
	S=> E(	2916	));
			
  U2964	: Soma_AMA3_1 PORT MAP(
	A=> C(	3028	),
	B=>E(	2855	),
	Cin=> Carry( 	2963	),
	Cout=> Carry( 	2964	),
	S=> E(	2917	));
			
  U2965	: Soma_AMA3_1 PORT MAP(
	A=> C(	3029	),
	B=>E(	2856	),
	Cin=> Carry( 	2964	),
	Cout=> Carry( 	2965	),
	S=> E(	2918	));
			
  U2966	: Soma_AMA3_1 PORT MAP(
	A=> C(	3030	),
	B=>E(	2857	),
	Cin=> Carry( 	2965	),
	Cout=> Carry( 	2966	),
	S=> E(	2919	));
			
  U2967	: Soma_AMA3_1 PORT MAP(
	A=> C(	3031	),
	B=>E(	2858	),
	Cin=> Carry( 	2966	),
	Cout=> Carry( 	2967	),
	S=> E(	2920	));
			
  U2968	: Soma_AMA3_1 PORT MAP(
	A=> C(	3032	),
	B=>E(	2859	),
	Cin=> Carry( 	2967	),
	Cout=> Carry( 	2968	),
	S=> E(	2921	));
			
  U2969	: Soma_AMA3_1 PORT MAP(
	A=> C(	3033	),
	B=>E(	2860	),
	Cin=> Carry( 	2968	),
	Cout=> Carry( 	2969	),
	S=> E(	2922	));
			
  U2970	: Soma_AMA3_1 PORT MAP(
	A=> C(	3034	),
	B=>E(	2861	),
	Cin=> Carry( 	2969	),
	Cout=> Carry( 	2970	),
	S=> E(	2923	));
			
  U2971	: Soma_AMA3_1 PORT MAP(
	A=> C(	3035	),
	B=>E(	2862	),
	Cin=> Carry( 	2970	),
	Cout=> Carry( 	2971	),
	S=> E(	2924	));
			
  U2972	: Soma_AMA3_1 PORT MAP(
	A=> C(	3036	),
	B=>E(	2863	),
	Cin=> Carry( 	2971	),
	Cout=> Carry( 	2972	),
	S=> E(	2925	));
			
  U2973	: Soma_AMA3_1 PORT MAP(
	A=> C(	3037	),
	B=>E(	2864	),
	Cin=> Carry( 	2972	),
	Cout=> Carry( 	2973	),
	S=> E(	2926	));
			
  U2974	: Soma_AMA3_1 PORT MAP(
	A=> C(	3038	),
	B=>E(	2865	),
	Cin=> Carry( 	2973	),
	Cout=> Carry( 	2974	),
	S=> E(	2927	));
			
  U2975	: Soma_AMA3_1 PORT MAP(
	A=> C(	3039	),
	B=>E(	2866	),
	Cin=> Carry( 	2974	),
	Cout=> Carry( 	2975	),
	S=> E(	2928	));
			
  U2976	: Soma_AMA3_1 PORT MAP(
	A=> C(	3040	),
	B=>E(	2867	),
	Cin=> Carry( 	2975	),
	Cout=> Carry( 	2976	),
	S=> E(	2929	));
			
  U2977	: Soma_AMA3_1 PORT MAP(
	A=> C(	3041	),
	B=>E(	2868	),
	Cin=> Carry( 	2976	),
	Cout=> Carry( 	2977	),
	S=> E(	2930	));
			
  U2978	: Soma_AMA3_1 PORT MAP(
	A=> C(	3042	),
	B=>E(	2869	),
	Cin=> Carry( 	2977	),
	Cout=> Carry( 	2978	),
	S=> E(	2931	));
			
  U2979	: Soma_AMA3_1 PORT MAP(
	A=> C(	3043	),
	B=>E(	2870	),
	Cin=> Carry( 	2978	),
	Cout=> Carry( 	2979	),
	S=> E(	2932	));
			
  U2980	: Soma_AMA3_1 PORT MAP(
	A=> C(	3044	),
	B=>E(	2871	),
	Cin=> Carry( 	2979	),
	Cout=> Carry( 	2980	),
	S=> E(	2933	));
			
  U2981	: Soma_AMA3_1 PORT MAP(
	A=> C(	3045	),
	B=>E(	2872	),
	Cin=> Carry( 	2980	),
	Cout=> Carry( 	2981	),
	S=> E(	2934	));
			
  U2982	: Soma_AMA3_1 PORT MAP(
	A=> C(	3046	),
	B=>E(	2873	),
	Cin=> Carry( 	2981	),
	Cout=> Carry( 	2982	),
	S=> E(	2935	));
			
  U2983	: Soma_AMA3_1 PORT MAP(
	A=> C(	3047	),
	B=>E(	2874	),
	Cin=> Carry( 	2982	),
	Cout=> Carry( 	2983	),
	S=> E(	2936	));
			
  U2984	: Soma_AMA3_1 PORT MAP(
	A=> C(	3048	),
	B=>E(	2875	),
	Cin=> Carry( 	2983	),
	Cout=> Carry( 	2984	),
	S=> E(	2937	));
			
  U2985	: Soma_AMA3_1 PORT MAP(
	A=> C(	3049	),
	B=>E(	2876	),
	Cin=> Carry( 	2984	),
	Cout=> Carry( 	2985	),
	S=> E(	2938	));
			
  U2986	: Soma_AMA3_1 PORT MAP(
	A=> C(	3050	),
	B=>E(	2877	),
	Cin=> Carry( 	2985	),
	Cout=> Carry( 	2986	),
	S=> E(	2939	));
			
  U2987	: Soma_AMA3_1 PORT MAP(
	A=> C(	3051	),
	B=>E(	2878	),
	Cin=> Carry( 	2986	),
	Cout=> Carry( 	2987	),
	S=> E(	2940	));
			
  U2988	: Soma_AMA3_1 PORT MAP(
	A=> C(	3052	),
	B=>E(	2879	),
	Cin=> Carry( 	2987	),
	Cout=> Carry( 	2988	),
	S=> E(	2941	));
			
  U2989	: Soma_AMA3_1 PORT MAP(
	A=> C(	3053	),
	B=>E(	2880	),
	Cin=> Carry( 	2988	),
	Cout=> Carry( 	2989	),
	S=> E(	2942	));
			
  U2990	: Soma_AMA3_1 PORT MAP(
	A=> C(	3054	),
	B=>E(	2881	),
	Cin=> Carry( 	2989	),
	Cout=> Carry( 	2990	),
	S=> E(	2943	));
			
  U2991	: Soma_AMA3_1 PORT MAP(
	A=> C(	3055	),
	B=>E(	2882	),
	Cin=> Carry( 	2990	),
	Cout=> Carry( 	2991	),
	S=> E(	2944	));
			
  U2992	: Soma_AMA3_1 PORT MAP(
	A=> C(	3056	),
	B=>E(	2883	),
	Cin=> Carry( 	2991	),
	Cout=> Carry( 	2992	),
	S=> E(	2945	));
			
  U2993	: Soma_AMA3_1 PORT MAP(
	A=> C(	3057	),
	B=>E(	2884	),
	Cin=> Carry( 	2992	),
	Cout=> Carry( 	2993	),
	S=> E(	2946	));
			
  U2994	: Soma_AMA3_1 PORT MAP(
	A=> C(	3058	),
	B=>E(	2885	),
	Cin=> Carry( 	2993	),
	Cout=> Carry( 	2994	),
	S=> E(	2947	));
			
  U2995	: Soma_AMA3_1 PORT MAP(
	A=> C(	3059	),
	B=>E(	2886	),
	Cin=> Carry( 	2994	),
	Cout=> Carry( 	2995	),
	S=> E(	2948	));
			
  U2996	: Soma_AMA3_1 PORT MAP(
	A=> C(	3060	),
	B=>E(	2887	),
	Cin=> Carry( 	2995	),
	Cout=> Carry( 	2996	),
	S=> E(	2949	));
			
  U2997	: Soma_AMA3_1 PORT MAP(
	A=> C(	3061	),
	B=>E(	2888	),
	Cin=> Carry( 	2996	),
	Cout=> Carry( 	2997	),
	S=> E(	2950	));
			
  U2998	: Soma_AMA3_1 PORT MAP(
	A=> C(	3062	),
	B=>E(	2889	),
	Cin=> Carry( 	2997	),
	Cout=> Carry( 	2998	),
	S=> E(	2951	));
			
  U2999	: Soma_AMA3_1 PORT MAP(
	A=> C(	3063	),
	B=>E(	2890	),
	Cin=> Carry( 	2998	),
	Cout=> Carry( 	2999	),
	S=> E(	2952	));
			
  U3000	: Soma_AMA3_1 PORT MAP(
	A=> C(	3064	),
	B=>E(	2891	),
	Cin=> Carry( 	2999	),
	Cout=> Carry( 	3000	),
	S=> E(	2953	));
			
  U3001	: Soma_AMA3_1 PORT MAP(
	A=> C(	3065	),
	B=>E(	2892	),
	Cin=> Carry( 	3000	),
	Cout=> Carry( 	3001	),
	S=> E(	2954	));
			
  U3002	: Soma_AMA3_1 PORT MAP(
	A=> C(	3066	),
	B=>E(	2893	),
	Cin=> Carry( 	3001	),
	Cout=> Carry( 	3002	),
	S=> E(	2955	));
			
  U3003	: Soma_AMA3_1 PORT MAP(
	A=> C(	3067	),
	B=>E(	2894	),
	Cin=> Carry( 	3002	),
	Cout=> Carry( 	3003	),
	S=> E(	2956	));
			
  U3004	: Soma_AMA3_1 PORT MAP(
	A=> C(	3068	),
	B=>E(	2895	),
	Cin=> Carry( 	3003	),
	Cout=> Carry( 	3004	),
	S=> E(	2957	));
			
  U3005	: Soma_AMA3_1 PORT MAP(
	A=> C(	3069	),
	B=>E(	2896	),
	Cin=> Carry( 	3004	),
	Cout=> Carry( 	3005	),
	S=> E(	2958	));
			
  U3006	: Soma_AMA3_1 PORT MAP(
	A=> C(	3070	),
	B=>E(	2897	),
	Cin=> Carry( 	3005	),
	Cout=> Carry( 	3006	),
	S=> E(	2959	));
			
  U3007	: Soma_AMA3_1 PORT MAP(
	A=> C(	3071	),
	B=>Carry(	2943	),
	Cin=> Carry( 	3006	),
	Cout=> Carry( 	3007	),
	S=> E(	2960	));

			
  U3008	: Soma_AMA3_1 PORT MAP(
	A=> C(	3072	),
	B=>E(	2898	),
	Cin=> '0'	,
	Cout=> Carry( 	3008	),
	S=> R(	48	));
			
  U3009	: Soma_AMA3_1 PORT MAP(
	A=> C(	3073	),
	B=>E(	2899	),
	Cin=> Carry( 	3008	),
	Cout=> Carry( 	3009	),
	S=> E(	2961	));
			
  U3010	: Soma_AMA3_1 PORT MAP(
	A=> C(	3074	),
	B=>E(	2900	),
	Cin=> Carry( 	3009	),
	Cout=> Carry( 	3010	),
	S=> E(	2962	));
			
  U3011	: Soma_AMA3_1 PORT MAP(
	A=> C(	3075	),
	B=>E(	2901	),
	Cin=> Carry( 	3010	),
	Cout=> Carry( 	3011	),
	S=> E(	2963	));
			
  U3012	: Soma_AMA3_1 PORT MAP(
	A=> C(	3076	),
	B=>E(	2902	),
	Cin=> Carry( 	3011	),
	Cout=> Carry( 	3012	),
	S=> E(	2964	));
			
  U3013	: Soma_AMA3_1 PORT MAP(
	A=> C(	3077	),
	B=>E(	2903	),
	Cin=> Carry( 	3012	),
	Cout=> Carry( 	3013	),
	S=> E(	2965	));
			
  U3014	: Soma_AMA3_1 PORT MAP(
	A=> C(	3078	),
	B=>E(	2904	),
	Cin=> Carry( 	3013	),
	Cout=> Carry( 	3014	),
	S=> E(	2966	));
			
  U3015	: Soma_AMA3_1 PORT MAP(
	A=> C(	3079	),
	B=>E(	2905	),
	Cin=> Carry( 	3014	),
	Cout=> Carry( 	3015	),
	S=> E(	2967	));
			
  U3016	: Soma_AMA3_1 PORT MAP(
	A=> C(	3080	),
	B=>E(	2906	),
	Cin=> Carry( 	3015	),
	Cout=> Carry( 	3016	),
	S=> E(	2968	));
			
  U3017	: Soma_AMA3_1 PORT MAP(
	A=> C(	3081	),
	B=>E(	2907	),
	Cin=> Carry( 	3016	),
	Cout=> Carry( 	3017	),
	S=> E(	2969	));
			
  U3018	: Soma_AMA3_1 PORT MAP(
	A=> C(	3082	),
	B=>E(	2908	),
	Cin=> Carry( 	3017	),
	Cout=> Carry( 	3018	),
	S=> E(	2970	));
			
  U3019	: Soma_AMA3_1 PORT MAP(
	A=> C(	3083	),
	B=>E(	2909	),
	Cin=> Carry( 	3018	),
	Cout=> Carry( 	3019	),
	S=> E(	2971	));
			
  U3020	: Soma_AMA3_1 PORT MAP(
	A=> C(	3084	),
	B=>E(	2910	),
	Cin=> Carry( 	3019	),
	Cout=> Carry( 	3020	),
	S=> E(	2972	));
			
  U3021	: Soma_AMA3_1 PORT MAP(
	A=> C(	3085	),
	B=>E(	2911	),
	Cin=> Carry( 	3020	),
	Cout=> Carry( 	3021	),
	S=> E(	2973	));
			
  U3022	: Soma_AMA3_1 PORT MAP(
	A=> C(	3086	),
	B=>E(	2912	),
	Cin=> Carry( 	3021	),
	Cout=> Carry( 	3022	),
	S=> E(	2974	));
			
  U3023	: Soma_AMA3_1 PORT MAP(
	A=> C(	3087	),
	B=>E(	2913	),
	Cin=> Carry( 	3022	),
	Cout=> Carry( 	3023	),
	S=> E(	2975	));
			
  U3024	: Soma_AMA3_1 PORT MAP(
	A=> C(	3088	),
	B=>E(	2914	),
	Cin=> Carry( 	3023	),
	Cout=> Carry( 	3024	),
	S=> E(	2976	));
			
  U3025	: Soma_AMA3_1 PORT MAP(
	A=> C(	3089	),
	B=>E(	2915	),
	Cin=> Carry( 	3024	),
	Cout=> Carry( 	3025	),
	S=> E(	2977	));
			
  U3026	: Soma_AMA3_1 PORT MAP(
	A=> C(	3090	),
	B=>E(	2916	),
	Cin=> Carry( 	3025	),
	Cout=> Carry( 	3026	),
	S=> E(	2978	));
			
  U3027	: Soma_AMA3_1 PORT MAP(
	A=> C(	3091	),
	B=>E(	2917	),
	Cin=> Carry( 	3026	),
	Cout=> Carry( 	3027	),
	S=> E(	2979	));
			
  U3028	: Soma_AMA3_1 PORT MAP(
	A=> C(	3092	),
	B=>E(	2918	),
	Cin=> Carry( 	3027	),
	Cout=> Carry( 	3028	),
	S=> E(	2980	));
			
  U3029	: Soma_AMA3_1 PORT MAP(
	A=> C(	3093	),
	B=>E(	2919	),
	Cin=> Carry( 	3028	),
	Cout=> Carry( 	3029	),
	S=> E(	2981	));
			
  U3030	: Soma_AMA3_1 PORT MAP(
	A=> C(	3094	),
	B=>E(	2920	),
	Cin=> Carry( 	3029	),
	Cout=> Carry( 	3030	),
	S=> E(	2982	));
			
  U3031	: Soma_AMA3_1 PORT MAP(
	A=> C(	3095	),
	B=>E(	2921	),
	Cin=> Carry( 	3030	),
	Cout=> Carry( 	3031	),
	S=> E(	2983	));
			
  U3032	: Soma_AMA3_1 PORT MAP(
	A=> C(	3096	),
	B=>E(	2922	),
	Cin=> Carry( 	3031	),
	Cout=> Carry( 	3032	),
	S=> E(	2984	));
			
  U3033	: Soma_AMA3_1 PORT MAP(
	A=> C(	3097	),
	B=>E(	2923	),
	Cin=> Carry( 	3032	),
	Cout=> Carry( 	3033	),
	S=> E(	2985	));
			
  U3034	: Soma_AMA3_1 PORT MAP(
	A=> C(	3098	),
	B=>E(	2924	),
	Cin=> Carry( 	3033	),
	Cout=> Carry( 	3034	),
	S=> E(	2986	));
			
  U3035	: Soma_AMA3_1 PORT MAP(
	A=> C(	3099	),
	B=>E(	2925	),
	Cin=> Carry( 	3034	),
	Cout=> Carry( 	3035	),
	S=> E(	2987	));
			
  U3036	: Soma_AMA3_1 PORT MAP(
	A=> C(	3100	),
	B=>E(	2926	),
	Cin=> Carry( 	3035	),
	Cout=> Carry( 	3036	),
	S=> E(	2988	));
			
  U3037	: Soma_AMA3_1 PORT MAP(
	A=> C(	3101	),
	B=>E(	2927	),
	Cin=> Carry( 	3036	),
	Cout=> Carry( 	3037	),
	S=> E(	2989	));
			
  U3038	: Soma_AMA3_1 PORT MAP(
	A=> C(	3102	),
	B=>E(	2928	),
	Cin=> Carry( 	3037	),
	Cout=> Carry( 	3038	),
	S=> E(	2990	));
			
  U3039	: Soma_AMA3_1 PORT MAP(
	A=> C(	3103	),
	B=>E(	2929	),
	Cin=> Carry( 	3038	),
	Cout=> Carry( 	3039	),
	S=> E(	2991	));
			
  U3040	: Soma_AMA3_1 PORT MAP(
	A=> C(	3104	),
	B=>E(	2930	),
	Cin=> Carry( 	3039	),
	Cout=> Carry( 	3040	),
	S=> E(	2992	));
			
  U3041	: Soma_AMA3_1 PORT MAP(
	A=> C(	3105	),
	B=>E(	2931	),
	Cin=> Carry( 	3040	),
	Cout=> Carry( 	3041	),
	S=> E(	2993	));
			
  U3042	: Soma_AMA3_1 PORT MAP(
	A=> C(	3106	),
	B=>E(	2932	),
	Cin=> Carry( 	3041	),
	Cout=> Carry( 	3042	),
	S=> E(	2994	));
			
  U3043	: Soma_AMA3_1 PORT MAP(
	A=> C(	3107	),
	B=>E(	2933	),
	Cin=> Carry( 	3042	),
	Cout=> Carry( 	3043	),
	S=> E(	2995	));
			
  U3044	: Soma_AMA3_1 PORT MAP(
	A=> C(	3108	),
	B=>E(	2934	),
	Cin=> Carry( 	3043	),
	Cout=> Carry( 	3044	),
	S=> E(	2996	));
			
  U3045	: Soma_AMA3_1 PORT MAP(
	A=> C(	3109	),
	B=>E(	2935	),
	Cin=> Carry( 	3044	),
	Cout=> Carry( 	3045	),
	S=> E(	2997	));
			
  U3046	: Soma_AMA3_1 PORT MAP(
	A=> C(	3110	),
	B=>E(	2936	),
	Cin=> Carry( 	3045	),
	Cout=> Carry( 	3046	),
	S=> E(	2998	));
			
  U3047	: Soma_AMA3_1 PORT MAP(
	A=> C(	3111	),
	B=>E(	2937	),
	Cin=> Carry( 	3046	),
	Cout=> Carry( 	3047	),
	S=> E(	2999	));
			
  U3048	: Soma_AMA3_1 PORT MAP(
	A=> C(	3112	),
	B=>E(	2938	),
	Cin=> Carry( 	3047	),
	Cout=> Carry( 	3048	),
	S=> E(	3000	));
			
  U3049	: Soma_AMA3_1 PORT MAP(
	A=> C(	3113	),
	B=>E(	2939	),
	Cin=> Carry( 	3048	),
	Cout=> Carry( 	3049	),
	S=> E(	3001	));
			
  U3050	: Soma_AMA3_1 PORT MAP(
	A=> C(	3114	),
	B=>E(	2940	),
	Cin=> Carry( 	3049	),
	Cout=> Carry( 	3050	),
	S=> E(	3002	));
			
  U3051	: Soma_AMA3_1 PORT MAP(
	A=> C(	3115	),
	B=>E(	2941	),
	Cin=> Carry( 	3050	),
	Cout=> Carry( 	3051	),
	S=> E(	3003	));
			
  U3052	: Soma_AMA3_1 PORT MAP(
	A=> C(	3116	),
	B=>E(	2942	),
	Cin=> Carry( 	3051	),
	Cout=> Carry( 	3052	),
	S=> E(	3004	));
			
  U3053	: Soma_AMA3_1 PORT MAP(
	A=> C(	3117	),
	B=>E(	2943	),
	Cin=> Carry( 	3052	),
	Cout=> Carry( 	3053	),
	S=> E(	3005	));
			
  U3054	: Soma_AMA3_1 PORT MAP(
	A=> C(	3118	),
	B=>E(	2944	),
	Cin=> Carry( 	3053	),
	Cout=> Carry( 	3054	),
	S=> E(	3006	));
			
  U3055	: Soma_AMA3_1 PORT MAP(
	A=> C(	3119	),
	B=>E(	2945	),
	Cin=> Carry( 	3054	),
	Cout=> Carry( 	3055	),
	S=> E(	3007	));
			
  U3056	: Soma_AMA3_1 PORT MAP(
	A=> C(	3120	),
	B=>E(	2946	),
	Cin=> Carry( 	3055	),
	Cout=> Carry( 	3056	),
	S=> E(	3008	));
			
  U3057	: Soma_AMA3_1 PORT MAP(
	A=> C(	3121	),
	B=>E(	2947	),
	Cin=> Carry( 	3056	),
	Cout=> Carry( 	3057	),
	S=> E(	3009	));
			
  U3058	: Soma_AMA3_1 PORT MAP(
	A=> C(	3122	),
	B=>E(	2948	),
	Cin=> Carry( 	3057	),
	Cout=> Carry( 	3058	),
	S=> E(	3010	));
			
  U3059	: Soma_AMA3_1 PORT MAP(
	A=> C(	3123	),
	B=>E(	2949	),
	Cin=> Carry( 	3058	),
	Cout=> Carry( 	3059	),
	S=> E(	3011	));
			
  U3060	: Soma_AMA3_1 PORT MAP(
	A=> C(	3124	),
	B=>E(	2950	),
	Cin=> Carry( 	3059	),
	Cout=> Carry( 	3060	),
	S=> E(	3012	));
			
  U3061	: Soma_AMA3_1 PORT MAP(
	A=> C(	3125	),
	B=>E(	2951	),
	Cin=> Carry( 	3060	),
	Cout=> Carry( 	3061	),
	S=> E(	3013	));
			
  U3062	: Soma_AMA3_1 PORT MAP(
	A=> C(	3126	),
	B=>E(	2952	),
	Cin=> Carry( 	3061	),
	Cout=> Carry( 	3062	),
	S=> E(	3014	));
			
  U3063	: Soma_AMA3_1 PORT MAP(
	A=> C(	3127	),
	B=>E(	2953	),
	Cin=> Carry( 	3062	),
	Cout=> Carry( 	3063	),
	S=> E(	3015	));
			
  U3064	: Soma_AMA3_1 PORT MAP(
	A=> C(	3128	),
	B=>E(	2954	),
	Cin=> Carry( 	3063	),
	Cout=> Carry( 	3064	),
	S=> E(	3016	));
			
  U3065	: Soma_AMA3_1 PORT MAP(
	A=> C(	3129	),
	B=>E(	2955	),
	Cin=> Carry( 	3064	),
	Cout=> Carry( 	3065	),
	S=> E(	3017	));
			
  U3066	: Soma_AMA3_1 PORT MAP(
	A=> C(	3130	),
	B=>E(	2956	),
	Cin=> Carry( 	3065	),
	Cout=> Carry( 	3066	),
	S=> E(	3018	));
			
  U3067	: Soma_AMA3_1 PORT MAP(
	A=> C(	3131	),
	B=>E(	2957	),
	Cin=> Carry( 	3066	),
	Cout=> Carry( 	3067	),
	S=> E(	3019	));
			
  U3068	: Soma_AMA3_1 PORT MAP(
	A=> C(	3132	),
	B=>E(	2958	),
	Cin=> Carry( 	3067	),
	Cout=> Carry( 	3068	),
	S=> E(	3020	));
			
  U3069	: Soma_AMA3_1 PORT MAP(
	A=> C(	3133	),
	B=>E(	2959	),
	Cin=> Carry( 	3068	),
	Cout=> Carry( 	3069	),
	S=> E(	3021	));
			
  U3070	: Soma_AMA3_1 PORT MAP(
	A=> C(	3134	),
	B=>E(	2960	),
	Cin=> Carry( 	3069	),
	Cout=> Carry( 	3070	),
	S=> E(	3022	));
			
  U3071	: Soma_AMA3_1 PORT MAP(
	A=> C(	3135	),
	B=>Carry(	3007	),
	Cin=> Carry( 	3070	),
	Cout=> Carry( 	3071	),
	S=> E(	3023	));

			
  U3072	: Soma_AMA3_1 PORT MAP(
	A=> C(	3136	),
	B=>E(	2961	),
	Cin=> '0'	,
	Cout=> Carry( 	3072	),
	S=> R(	49	));
			
  U3073	: Soma_AMA3_1 PORT MAP(
	A=> C(	3137	),
	B=>E(	2962	),
	Cin=> Carry( 	3072	),
	Cout=> Carry( 	3073	),
	S=> E(	3024	));
			
  U3074	: Soma_AMA3_1 PORT MAP(
	A=> C(	3138	),
	B=>E(	2963	),
	Cin=> Carry( 	3073	),
	Cout=> Carry( 	3074	),
	S=> E(	3025	));
			
  U3075	: Soma_AMA3_1 PORT MAP(
	A=> C(	3139	),
	B=>E(	2964	),
	Cin=> Carry( 	3074	),
	Cout=> Carry( 	3075	),
	S=> E(	3026	));
			
  U3076	: Soma_AMA3_1 PORT MAP(
	A=> C(	3140	),
	B=>E(	2965	),
	Cin=> Carry( 	3075	),
	Cout=> Carry( 	3076	),
	S=> E(	3027	));
			
  U3077	: Soma_AMA3_1 PORT MAP(
	A=> C(	3141	),
	B=>E(	2966	),
	Cin=> Carry( 	3076	),
	Cout=> Carry( 	3077	),
	S=> E(	3028	));
			
  U3078	: Soma_AMA3_1 PORT MAP(
	A=> C(	3142	),
	B=>E(	2967	),
	Cin=> Carry( 	3077	),
	Cout=> Carry( 	3078	),
	S=> E(	3029	));
			
  U3079	: Soma_AMA3_1 PORT MAP(
	A=> C(	3143	),
	B=>E(	2968	),
	Cin=> Carry( 	3078	),
	Cout=> Carry( 	3079	),
	S=> E(	3030	));
			
  U3080	: Soma_AMA3_1 PORT MAP(
	A=> C(	3144	),
	B=>E(	2969	),
	Cin=> Carry( 	3079	),
	Cout=> Carry( 	3080	),
	S=> E(	3031	));
			
  U3081	: Soma_AMA3_1 PORT MAP(
	A=> C(	3145	),
	B=>E(	2970	),
	Cin=> Carry( 	3080	),
	Cout=> Carry( 	3081	),
	S=> E(	3032	));
			
  U3082	: Soma_AMA3_1 PORT MAP(
	A=> C(	3146	),
	B=>E(	2971	),
	Cin=> Carry( 	3081	),
	Cout=> Carry( 	3082	),
	S=> E(	3033	));
			
  U3083	: Soma_AMA3_1 PORT MAP(
	A=> C(	3147	),
	B=>E(	2972	),
	Cin=> Carry( 	3082	),
	Cout=> Carry( 	3083	),
	S=> E(	3034	));
			
  U3084	: Soma_AMA3_1 PORT MAP(
	A=> C(	3148	),
	B=>E(	2973	),
	Cin=> Carry( 	3083	),
	Cout=> Carry( 	3084	),
	S=> E(	3035	));
			
  U3085	: Soma_AMA3_1 PORT MAP(
	A=> C(	3149	),
	B=>E(	2974	),
	Cin=> Carry( 	3084	),
	Cout=> Carry( 	3085	),
	S=> E(	3036	));
			
  U3086	: Soma_AMA3_1 PORT MAP(
	A=> C(	3150	),
	B=>E(	2975	),
	Cin=> Carry( 	3085	),
	Cout=> Carry( 	3086	),
	S=> E(	3037	));
			
  U3087	: Soma_AMA3_1 PORT MAP(
	A=> C(	3151	),
	B=>E(	2976	),
	Cin=> Carry( 	3086	),
	Cout=> Carry( 	3087	),
	S=> E(	3038	));
			
  U3088	: Soma_AMA3_1 PORT MAP(
	A=> C(	3152	),
	B=>E(	2977	),
	Cin=> Carry( 	3087	),
	Cout=> Carry( 	3088	),
	S=> E(	3039	));
			
  U3089	: Soma_AMA3_1 PORT MAP(
	A=> C(	3153	),
	B=>E(	2978	),
	Cin=> Carry( 	3088	),
	Cout=> Carry( 	3089	),
	S=> E(	3040	));
			
  U3090	: Soma_AMA3_1 PORT MAP(
	A=> C(	3154	),
	B=>E(	2979	),
	Cin=> Carry( 	3089	),
	Cout=> Carry( 	3090	),
	S=> E(	3041	));
			
  U3091	: Soma_AMA3_1 PORT MAP(
	A=> C(	3155	),
	B=>E(	2980	),
	Cin=> Carry( 	3090	),
	Cout=> Carry( 	3091	),
	S=> E(	3042	));
			
  U3092	: Soma_AMA3_1 PORT MAP(
	A=> C(	3156	),
	B=>E(	2981	),
	Cin=> Carry( 	3091	),
	Cout=> Carry( 	3092	),
	S=> E(	3043	));
			
  U3093	: Soma_AMA3_1 PORT MAP(
	A=> C(	3157	),
	B=>E(	2982	),
	Cin=> Carry( 	3092	),
	Cout=> Carry( 	3093	),
	S=> E(	3044	));
			
  U3094	: Soma_AMA3_1 PORT MAP(
	A=> C(	3158	),
	B=>E(	2983	),
	Cin=> Carry( 	3093	),
	Cout=> Carry( 	3094	),
	S=> E(	3045	));
			
  U3095	: Soma_AMA3_1 PORT MAP(
	A=> C(	3159	),
	B=>E(	2984	),
	Cin=> Carry( 	3094	),
	Cout=> Carry( 	3095	),
	S=> E(	3046	));
			
  U3096	: Soma_AMA3_1 PORT MAP(
	A=> C(	3160	),
	B=>E(	2985	),
	Cin=> Carry( 	3095	),
	Cout=> Carry( 	3096	),
	S=> E(	3047	));
			
  U3097	: Soma_AMA3_1 PORT MAP(
	A=> C(	3161	),
	B=>E(	2986	),
	Cin=> Carry( 	3096	),
	Cout=> Carry( 	3097	),
	S=> E(	3048	));
			
  U3098	: Soma_AMA3_1 PORT MAP(
	A=> C(	3162	),
	B=>E(	2987	),
	Cin=> Carry( 	3097	),
	Cout=> Carry( 	3098	),
	S=> E(	3049	));
			
  U3099	: Soma_AMA3_1 PORT MAP(
	A=> C(	3163	),
	B=>E(	2988	),
	Cin=> Carry( 	3098	),
	Cout=> Carry( 	3099	),
	S=> E(	3050	));
			
  U3100	: Soma_AMA3_1 PORT MAP(
	A=> C(	3164	),
	B=>E(	2989	),
	Cin=> Carry( 	3099	),
	Cout=> Carry( 	3100	),
	S=> E(	3051	));
			
  U3101	: Soma_AMA3_1 PORT MAP(
	A=> C(	3165	),
	B=>E(	2990	),
	Cin=> Carry( 	3100	),
	Cout=> Carry( 	3101	),
	S=> E(	3052	));
			
  U3102	: Soma_AMA3_1 PORT MAP(
	A=> C(	3166	),
	B=>E(	2991	),
	Cin=> Carry( 	3101	),
	Cout=> Carry( 	3102	),
	S=> E(	3053	));
			
  U3103	: Soma_AMA3_1 PORT MAP(
	A=> C(	3167	),
	B=>E(	2992	),
	Cin=> Carry( 	3102	),
	Cout=> Carry( 	3103	),
	S=> E(	3054	));
			
  U3104	: Soma_AMA3_1 PORT MAP(
	A=> C(	3168	),
	B=>E(	2993	),
	Cin=> Carry( 	3103	),
	Cout=> Carry( 	3104	),
	S=> E(	3055	));
			
  U3105	: Soma_AMA3_1 PORT MAP(
	A=> C(	3169	),
	B=>E(	2994	),
	Cin=> Carry( 	3104	),
	Cout=> Carry( 	3105	),
	S=> E(	3056	));
			
  U3106	: Soma_AMA3_1 PORT MAP(
	A=> C(	3170	),
	B=>E(	2995	),
	Cin=> Carry( 	3105	),
	Cout=> Carry( 	3106	),
	S=> E(	3057	));
			
  U3107	: Soma_AMA3_1 PORT MAP(
	A=> C(	3171	),
	B=>E(	2996	),
	Cin=> Carry( 	3106	),
	Cout=> Carry( 	3107	),
	S=> E(	3058	));
			
  U3108	: Soma_AMA3_1 PORT MAP(
	A=> C(	3172	),
	B=>E(	2997	),
	Cin=> Carry( 	3107	),
	Cout=> Carry( 	3108	),
	S=> E(	3059	));
			
  U3109	: Soma_AMA3_1 PORT MAP(
	A=> C(	3173	),
	B=>E(	2998	),
	Cin=> Carry( 	3108	),
	Cout=> Carry( 	3109	),
	S=> E(	3060	));
			
  U3110	: Soma_AMA3_1 PORT MAP(
	A=> C(	3174	),
	B=>E(	2999	),
	Cin=> Carry( 	3109	),
	Cout=> Carry( 	3110	),
	S=> E(	3061	));
			
  U3111	: Soma_AMA3_1 PORT MAP(
	A=> C(	3175	),
	B=>E(	3000	),
	Cin=> Carry( 	3110	),
	Cout=> Carry( 	3111	),
	S=> E(	3062	));
			
  U3112	: Soma_AMA3_1 PORT MAP(
	A=> C(	3176	),
	B=>E(	3001	),
	Cin=> Carry( 	3111	),
	Cout=> Carry( 	3112	),
	S=> E(	3063	));
			
  U3113	: Soma_AMA3_1 PORT MAP(
	A=> C(	3177	),
	B=>E(	3002	),
	Cin=> Carry( 	3112	),
	Cout=> Carry( 	3113	),
	S=> E(	3064	));
			
  U3114	: Soma_AMA3_1 PORT MAP(
	A=> C(	3178	),
	B=>E(	3003	),
	Cin=> Carry( 	3113	),
	Cout=> Carry( 	3114	),
	S=> E(	3065	));
			
  U3115	: Soma_AMA3_1 PORT MAP(
	A=> C(	3179	),
	B=>E(	3004	),
	Cin=> Carry( 	3114	),
	Cout=> Carry( 	3115	),
	S=> E(	3066	));
			
  U3116	: Soma_AMA3_1 PORT MAP(
	A=> C(	3180	),
	B=>E(	3005	),
	Cin=> Carry( 	3115	),
	Cout=> Carry( 	3116	),
	S=> E(	3067	));
			
  U3117	: Soma_AMA3_1 PORT MAP(
	A=> C(	3181	),
	B=>E(	3006	),
	Cin=> Carry( 	3116	),
	Cout=> Carry( 	3117	),
	S=> E(	3068	));
			
  U3118	: Soma_AMA3_1 PORT MAP(
	A=> C(	3182	),
	B=>E(	3007	),
	Cin=> Carry( 	3117	),
	Cout=> Carry( 	3118	),
	S=> E(	3069	));
			
  U3119	: Soma_AMA3_1 PORT MAP(
	A=> C(	3183	),
	B=>E(	3008	),
	Cin=> Carry( 	3118	),
	Cout=> Carry( 	3119	),
	S=> E(	3070	));
			
  U3120	: Soma_AMA3_1 PORT MAP(
	A=> C(	3184	),
	B=>E(	3009	),
	Cin=> Carry( 	3119	),
	Cout=> Carry( 	3120	),
	S=> E(	3071	));
			
  U3121	: Soma_AMA3_1 PORT MAP(
	A=> C(	3185	),
	B=>E(	3010	),
	Cin=> Carry( 	3120	),
	Cout=> Carry( 	3121	),
	S=> E(	3072	));
			
  U3122	: Soma_AMA3_1 PORT MAP(
	A=> C(	3186	),
	B=>E(	3011	),
	Cin=> Carry( 	3121	),
	Cout=> Carry( 	3122	),
	S=> E(	3073	));
			
  U3123	: Soma_AMA3_1 PORT MAP(
	A=> C(	3187	),
	B=>E(	3012	),
	Cin=> Carry( 	3122	),
	Cout=> Carry( 	3123	),
	S=> E(	3074	));
			
  U3124	: Soma_AMA3_1 PORT MAP(
	A=> C(	3188	),
	B=>E(	3013	),
	Cin=> Carry( 	3123	),
	Cout=> Carry( 	3124	),
	S=> E(	3075	));
			
  U3125	: Soma_AMA3_1 PORT MAP(
	A=> C(	3189	),
	B=>E(	3014	),
	Cin=> Carry( 	3124	),
	Cout=> Carry( 	3125	),
	S=> E(	3076	));
			
  U3126	: Soma_AMA3_1 PORT MAP(
	A=> C(	3190	),
	B=>E(	3015	),
	Cin=> Carry( 	3125	),
	Cout=> Carry( 	3126	),
	S=> E(	3077	));
			
  U3127	: Soma_AMA3_1 PORT MAP(
	A=> C(	3191	),
	B=>E(	3016	),
	Cin=> Carry( 	3126	),
	Cout=> Carry( 	3127	),
	S=> E(	3078	));
			
  U3128	: Soma_AMA3_1 PORT MAP(
	A=> C(	3192	),
	B=>E(	3017	),
	Cin=> Carry( 	3127	),
	Cout=> Carry( 	3128	),
	S=> E(	3079	));
			
  U3129	: Soma_AMA3_1 PORT MAP(
	A=> C(	3193	),
	B=>E(	3018	),
	Cin=> Carry( 	3128	),
	Cout=> Carry( 	3129	),
	S=> E(	3080	));
			
  U3130	: Soma_AMA3_1 PORT MAP(
	A=> C(	3194	),
	B=>E(	3019	),
	Cin=> Carry( 	3129	),
	Cout=> Carry( 	3130	),
	S=> E(	3081	));
			
  U3131	: Soma_AMA3_1 PORT MAP(
	A=> C(	3195	),
	B=>E(	3020	),
	Cin=> Carry( 	3130	),
	Cout=> Carry( 	3131	),
	S=> E(	3082	));
			
  U3132	: Soma_AMA3_1 PORT MAP(
	A=> C(	3196	),
	B=>E(	3021	),
	Cin=> Carry( 	3131	),
	Cout=> Carry( 	3132	),
	S=> E(	3083	));
			
  U3133	: Soma_AMA3_1 PORT MAP(
	A=> C(	3197	),
	B=>E(	3022	),
	Cin=> Carry( 	3132	),
	Cout=> Carry( 	3133	),
	S=> E(	3084	));
			
  U3134	: Soma_AMA3_1 PORT MAP(
	A=> C(	3198	),
	B=>E(	3023	),
	Cin=> Carry( 	3133	),
	Cout=> Carry( 	3134	),
	S=> E(	3085	));
			
  U3135	: Soma_AMA3_1 PORT MAP(
	A=> C(	3199	),
	B=>Carry(	3071	),
	Cin=> Carry( 	3134	),
	Cout=> Carry( 	3135	),
	S=> E(	3086	));

			
  U3136	: Soma_AMA3_1 PORT MAP(
	A=> C(	3200	),
	B=>E(	3024	),
	Cin=> '0'	,
	Cout=> Carry( 	3136	),
	S=> R(	50	));
			
  U3137	: Soma_AMA3_1 PORT MAP(
	A=> C(	3201	),
	B=>E(	3025	),
	Cin=> Carry( 	3136	),
	Cout=> Carry( 	3137	),
	S=> E(	3087	));
			
  U3138	: Soma_AMA3_1 PORT MAP(
	A=> C(	3202	),
	B=>E(	3026	),
	Cin=> Carry( 	3137	),
	Cout=> Carry( 	3138	),
	S=> E(	3088	));
			
  U3139	: Soma_AMA3_1 PORT MAP(
	A=> C(	3203	),
	B=>E(	3027	),
	Cin=> Carry( 	3138	),
	Cout=> Carry( 	3139	),
	S=> E(	3089	));
			
  U3140	: Soma_AMA3_1 PORT MAP(
	A=> C(	3204	),
	B=>E(	3028	),
	Cin=> Carry( 	3139	),
	Cout=> Carry( 	3140	),
	S=> E(	3090	));
			
  U3141	: Soma_AMA3_1 PORT MAP(
	A=> C(	3205	),
	B=>E(	3029	),
	Cin=> Carry( 	3140	),
	Cout=> Carry( 	3141	),
	S=> E(	3091	));
			
  U3142	: Soma_AMA3_1 PORT MAP(
	A=> C(	3206	),
	B=>E(	3030	),
	Cin=> Carry( 	3141	),
	Cout=> Carry( 	3142	),
	S=> E(	3092	));
			
  U3143	: Soma_AMA3_1 PORT MAP(
	A=> C(	3207	),
	B=>E(	3031	),
	Cin=> Carry( 	3142	),
	Cout=> Carry( 	3143	),
	S=> E(	3093	));
			
  U3144	: Soma_AMA3_1 PORT MAP(
	A=> C(	3208	),
	B=>E(	3032	),
	Cin=> Carry( 	3143	),
	Cout=> Carry( 	3144	),
	S=> E(	3094	));
			
  U3145	: Soma_AMA3_1 PORT MAP(
	A=> C(	3209	),
	B=>E(	3033	),
	Cin=> Carry( 	3144	),
	Cout=> Carry( 	3145	),
	S=> E(	3095	));
			
  U3146	: Soma_AMA3_1 PORT MAP(
	A=> C(	3210	),
	B=>E(	3034	),
	Cin=> Carry( 	3145	),
	Cout=> Carry( 	3146	),
	S=> E(	3096	));
			
  U3147	: Soma_AMA3_1 PORT MAP(
	A=> C(	3211	),
	B=>E(	3035	),
	Cin=> Carry( 	3146	),
	Cout=> Carry( 	3147	),
	S=> E(	3097	));
			
  U3148	: Soma_AMA3_1 PORT MAP(
	A=> C(	3212	),
	B=>E(	3036	),
	Cin=> Carry( 	3147	),
	Cout=> Carry( 	3148	),
	S=> E(	3098	));
			
  U3149	: Soma_AMA3_1 PORT MAP(
	A=> C(	3213	),
	B=>E(	3037	),
	Cin=> Carry( 	3148	),
	Cout=> Carry( 	3149	),
	S=> E(	3099	));
			
  U3150	: Soma_AMA3_1 PORT MAP(
	A=> C(	3214	),
	B=>E(	3038	),
	Cin=> Carry( 	3149	),
	Cout=> Carry( 	3150	),
	S=> E(	3100	));
			
  U3151	: Soma_AMA3_1 PORT MAP(
	A=> C(	3215	),
	B=>E(	3039	),
	Cin=> Carry( 	3150	),
	Cout=> Carry( 	3151	),
	S=> E(	3101	));
			
  U3152	: Soma_AMA3_1 PORT MAP(
	A=> C(	3216	),
	B=>E(	3040	),
	Cin=> Carry( 	3151	),
	Cout=> Carry( 	3152	),
	S=> E(	3102	));
			
  U3153	: Soma_AMA3_1 PORT MAP(
	A=> C(	3217	),
	B=>E(	3041	),
	Cin=> Carry( 	3152	),
	Cout=> Carry( 	3153	),
	S=> E(	3103	));
			
  U3154	: Soma_AMA3_1 PORT MAP(
	A=> C(	3218	),
	B=>E(	3042	),
	Cin=> Carry( 	3153	),
	Cout=> Carry( 	3154	),
	S=> E(	3104	));
			
  U3155	: Soma_AMA3_1 PORT MAP(
	A=> C(	3219	),
	B=>E(	3043	),
	Cin=> Carry( 	3154	),
	Cout=> Carry( 	3155	),
	S=> E(	3105	));
			
  U3156	: Soma_AMA3_1 PORT MAP(
	A=> C(	3220	),
	B=>E(	3044	),
	Cin=> Carry( 	3155	),
	Cout=> Carry( 	3156	),
	S=> E(	3106	));
			
  U3157	: Soma_AMA3_1 PORT MAP(
	A=> C(	3221	),
	B=>E(	3045	),
	Cin=> Carry( 	3156	),
	Cout=> Carry( 	3157	),
	S=> E(	3107	));
			
  U3158	: Soma_AMA3_1 PORT MAP(
	A=> C(	3222	),
	B=>E(	3046	),
	Cin=> Carry( 	3157	),
	Cout=> Carry( 	3158	),
	S=> E(	3108	));
			
  U3159	: Soma_AMA3_1 PORT MAP(
	A=> C(	3223	),
	B=>E(	3047	),
	Cin=> Carry( 	3158	),
	Cout=> Carry( 	3159	),
	S=> E(	3109	));
			
  U3160	: Soma_AMA3_1 PORT MAP(
	A=> C(	3224	),
	B=>E(	3048	),
	Cin=> Carry( 	3159	),
	Cout=> Carry( 	3160	),
	S=> E(	3110	));
			
  U3161	: Soma_AMA3_1 PORT MAP(
	A=> C(	3225	),
	B=>E(	3049	),
	Cin=> Carry( 	3160	),
	Cout=> Carry( 	3161	),
	S=> E(	3111	));
			
  U3162	: Soma_AMA3_1 PORT MAP(
	A=> C(	3226	),
	B=>E(	3050	),
	Cin=> Carry( 	3161	),
	Cout=> Carry( 	3162	),
	S=> E(	3112	));
			
  U3163	: Soma_AMA3_1 PORT MAP(
	A=> C(	3227	),
	B=>E(	3051	),
	Cin=> Carry( 	3162	),
	Cout=> Carry( 	3163	),
	S=> E(	3113	));
			
  U3164	: Soma_AMA3_1 PORT MAP(
	A=> C(	3228	),
	B=>E(	3052	),
	Cin=> Carry( 	3163	),
	Cout=> Carry( 	3164	),
	S=> E(	3114	));
			
  U3165	: Soma_AMA3_1 PORT MAP(
	A=> C(	3229	),
	B=>E(	3053	),
	Cin=> Carry( 	3164	),
	Cout=> Carry( 	3165	),
	S=> E(	3115	));
			
  U3166	: Soma_AMA3_1 PORT MAP(
	A=> C(	3230	),
	B=>E(	3054	),
	Cin=> Carry( 	3165	),
	Cout=> Carry( 	3166	),
	S=> E(	3116	));
			
  U3167	: Soma_AMA3_1 PORT MAP(
	A=> C(	3231	),
	B=>E(	3055	),
	Cin=> Carry( 	3166	),
	Cout=> Carry( 	3167	),
	S=> E(	3117	));
			
  U3168	: Soma_AMA3_1 PORT MAP(
	A=> C(	3232	),
	B=>E(	3056	),
	Cin=> Carry( 	3167	),
	Cout=> Carry( 	3168	),
	S=> E(	3118	));
			
  U3169	: Soma_AMA3_1 PORT MAP(
	A=> C(	3233	),
	B=>E(	3057	),
	Cin=> Carry( 	3168	),
	Cout=> Carry( 	3169	),
	S=> E(	3119	));
			
  U3170	: Soma_AMA3_1 PORT MAP(
	A=> C(	3234	),
	B=>E(	3058	),
	Cin=> Carry( 	3169	),
	Cout=> Carry( 	3170	),
	S=> E(	3120	));
			
  U3171	: Soma_AMA3_1 PORT MAP(
	A=> C(	3235	),
	B=>E(	3059	),
	Cin=> Carry( 	3170	),
	Cout=> Carry( 	3171	),
	S=> E(	3121	));
			
  U3172	: Soma_AMA3_1 PORT MAP(
	A=> C(	3236	),
	B=>E(	3060	),
	Cin=> Carry( 	3171	),
	Cout=> Carry( 	3172	),
	S=> E(	3122	));
			
  U3173	: Soma_AMA3_1 PORT MAP(
	A=> C(	3237	),
	B=>E(	3061	),
	Cin=> Carry( 	3172	),
	Cout=> Carry( 	3173	),
	S=> E(	3123	));
			
  U3174	: Soma_AMA3_1 PORT MAP(
	A=> C(	3238	),
	B=>E(	3062	),
	Cin=> Carry( 	3173	),
	Cout=> Carry( 	3174	),
	S=> E(	3124	));
			
  U3175	: Soma_AMA3_1 PORT MAP(
	A=> C(	3239	),
	B=>E(	3063	),
	Cin=> Carry( 	3174	),
	Cout=> Carry( 	3175	),
	S=> E(	3125	));
			
  U3176	: Soma_AMA3_1 PORT MAP(
	A=> C(	3240	),
	B=>E(	3064	),
	Cin=> Carry( 	3175	),
	Cout=> Carry( 	3176	),
	S=> E(	3126	));
			
  U3177	: Soma_AMA3_1 PORT MAP(
	A=> C(	3241	),
	B=>E(	3065	),
	Cin=> Carry( 	3176	),
	Cout=> Carry( 	3177	),
	S=> E(	3127	));
			
  U3178	: Soma_AMA3_1 PORT MAP(
	A=> C(	3242	),
	B=>E(	3066	),
	Cin=> Carry( 	3177	),
	Cout=> Carry( 	3178	),
	S=> E(	3128	));
			
  U3179	: Soma_AMA3_1 PORT MAP(
	A=> C(	3243	),
	B=>E(	3067	),
	Cin=> Carry( 	3178	),
	Cout=> Carry( 	3179	),
	S=> E(	3129	));
			
  U3180	: Soma_AMA3_1 PORT MAP(
	A=> C(	3244	),
	B=>E(	3068	),
	Cin=> Carry( 	3179	),
	Cout=> Carry( 	3180	),
	S=> E(	3130	));
			
  U3181	: Soma_AMA3_1 PORT MAP(
	A=> C(	3245	),
	B=>E(	3069	),
	Cin=> Carry( 	3180	),
	Cout=> Carry( 	3181	),
	S=> E(	3131	));
			
  U3182	: Soma_AMA3_1 PORT MAP(
	A=> C(	3246	),
	B=>E(	3070	),
	Cin=> Carry( 	3181	),
	Cout=> Carry( 	3182	),
	S=> E(	3132	));
			
  U3183	: Soma_AMA3_1 PORT MAP(
	A=> C(	3247	),
	B=>E(	3071	),
	Cin=> Carry( 	3182	),
	Cout=> Carry( 	3183	),
	S=> E(	3133	));
			
  U3184	: Soma_AMA3_1 PORT MAP(
	A=> C(	3248	),
	B=>E(	3072	),
	Cin=> Carry( 	3183	),
	Cout=> Carry( 	3184	),
	S=> E(	3134	));
			
  U3185	: Soma_AMA3_1 PORT MAP(
	A=> C(	3249	),
	B=>E(	3073	),
	Cin=> Carry( 	3184	),
	Cout=> Carry( 	3185	),
	S=> E(	3135	));
			
  U3186	: Soma_AMA3_1 PORT MAP(
	A=> C(	3250	),
	B=>E(	3074	),
	Cin=> Carry( 	3185	),
	Cout=> Carry( 	3186	),
	S=> E(	3136	));
			
  U3187	: Soma_AMA3_1 PORT MAP(
	A=> C(	3251	),
	B=>E(	3075	),
	Cin=> Carry( 	3186	),
	Cout=> Carry( 	3187	),
	S=> E(	3137	));
			
  U3188	: Soma_AMA3_1 PORT MAP(
	A=> C(	3252	),
	B=>E(	3076	),
	Cin=> Carry( 	3187	),
	Cout=> Carry( 	3188	),
	S=> E(	3138	));
			
  U3189	: Soma_AMA3_1 PORT MAP(
	A=> C(	3253	),
	B=>E(	3077	),
	Cin=> Carry( 	3188	),
	Cout=> Carry( 	3189	),
	S=> E(	3139	));
			
  U3190	: Soma_AMA3_1 PORT MAP(
	A=> C(	3254	),
	B=>E(	3078	),
	Cin=> Carry( 	3189	),
	Cout=> Carry( 	3190	),
	S=> E(	3140	));
			
  U3191	: Soma_AMA3_1 PORT MAP(
	A=> C(	3255	),
	B=>E(	3079	),
	Cin=> Carry( 	3190	),
	Cout=> Carry( 	3191	),
	S=> E(	3141	));
			
  U3192	: Soma_AMA3_1 PORT MAP(
	A=> C(	3256	),
	B=>E(	3080	),
	Cin=> Carry( 	3191	),
	Cout=> Carry( 	3192	),
	S=> E(	3142	));
			
  U3193	: Soma_AMA3_1 PORT MAP(
	A=> C(	3257	),
	B=>E(	3081	),
	Cin=> Carry( 	3192	),
	Cout=> Carry( 	3193	),
	S=> E(	3143	));
			
  U3194	: Soma_AMA3_1 PORT MAP(
	A=> C(	3258	),
	B=>E(	3082	),
	Cin=> Carry( 	3193	),
	Cout=> Carry( 	3194	),
	S=> E(	3144	));
			
  U3195	: Soma_AMA3_1 PORT MAP(
	A=> C(	3259	),
	B=>E(	3083	),
	Cin=> Carry( 	3194	),
	Cout=> Carry( 	3195	),
	S=> E(	3145	));
			
  U3196	: Soma_AMA3_1 PORT MAP(
	A=> C(	3260	),
	B=>E(	3084	),
	Cin=> Carry( 	3195	),
	Cout=> Carry( 	3196	),
	S=> E(	3146	));
			
  U3197	: Soma_AMA3_1 PORT MAP(
	A=> C(	3261	),
	B=>E(	3085	),
	Cin=> Carry( 	3196	),
	Cout=> Carry( 	3197	),
	S=> E(	3147	));
			
  U3198	: Soma_AMA3_1 PORT MAP(
	A=> C(	3262	),
	B=>E(	3086	),
	Cin=> Carry( 	3197	),
	Cout=> Carry( 	3198	),
	S=> E(	3148	));
			
  U3199	: Soma_AMA3_1 PORT MAP(
	A=> C(	3263	),
	B=>Carry(	3135	),
	Cin=> Carry( 	3198	),
	Cout=> Carry( 	3199	),
	S=> E(	3149	));

			
  U3200	: Soma_AMA3_1 PORT MAP(
	A=> C(	3264	),
	B=>E(	3087	),
	Cin=> '0'	,
	Cout=> Carry( 	3200	),
	S=> R(	51	));
			
  U3201	: Soma_AMA3_1 PORT MAP(
	A=> C(	3265	),
	B=>E(	3088	),
	Cin=> Carry( 	3200	),
	Cout=> Carry( 	3201	),
	S=> E(	3150	));
			
  U3202	: Soma_AMA3_1 PORT MAP(
	A=> C(	3266	),
	B=>E(	3089	),
	Cin=> Carry( 	3201	),
	Cout=> Carry( 	3202	),
	S=> E(	3151	));
			
  U3203	: Soma_AMA3_1 PORT MAP(
	A=> C(	3267	),
	B=>E(	3090	),
	Cin=> Carry( 	3202	),
	Cout=> Carry( 	3203	),
	S=> E(	3152	));
			
  U3204	: Soma_AMA3_1 PORT MAP(
	A=> C(	3268	),
	B=>E(	3091	),
	Cin=> Carry( 	3203	),
	Cout=> Carry( 	3204	),
	S=> E(	3153	));
			
  U3205	: Soma_AMA3_1 PORT MAP(
	A=> C(	3269	),
	B=>E(	3092	),
	Cin=> Carry( 	3204	),
	Cout=> Carry( 	3205	),
	S=> E(	3154	));
			
  U3206	: Soma_AMA3_1 PORT MAP(
	A=> C(	3270	),
	B=>E(	3093	),
	Cin=> Carry( 	3205	),
	Cout=> Carry( 	3206	),
	S=> E(	3155	));
			
  U3207	: Soma_AMA3_1 PORT MAP(
	A=> C(	3271	),
	B=>E(	3094	),
	Cin=> Carry( 	3206	),
	Cout=> Carry( 	3207	),
	S=> E(	3156	));
			
  U3208	: Soma_AMA3_1 PORT MAP(
	A=> C(	3272	),
	B=>E(	3095	),
	Cin=> Carry( 	3207	),
	Cout=> Carry( 	3208	),
	S=> E(	3157	));
			
  U3209	: Soma_AMA3_1 PORT MAP(
	A=> C(	3273	),
	B=>E(	3096	),
	Cin=> Carry( 	3208	),
	Cout=> Carry( 	3209	),
	S=> E(	3158	));
			
  U3210	: Soma_AMA3_1 PORT MAP(
	A=> C(	3274	),
	B=>E(	3097	),
	Cin=> Carry( 	3209	),
	Cout=> Carry( 	3210	),
	S=> E(	3159	));
			
  U3211	: Soma_AMA3_1 PORT MAP(
	A=> C(	3275	),
	B=>E(	3098	),
	Cin=> Carry( 	3210	),
	Cout=> Carry( 	3211	),
	S=> E(	3160	));
			
  U3212	: Soma_AMA3_1 PORT MAP(
	A=> C(	3276	),
	B=>E(	3099	),
	Cin=> Carry( 	3211	),
	Cout=> Carry( 	3212	),
	S=> E(	3161	));
			
  U3213	: Soma_AMA3_1 PORT MAP(
	A=> C(	3277	),
	B=>E(	3100	),
	Cin=> Carry( 	3212	),
	Cout=> Carry( 	3213	),
	S=> E(	3162	));
			
  U3214	: Soma_AMA3_1 PORT MAP(
	A=> C(	3278	),
	B=>E(	3101	),
	Cin=> Carry( 	3213	),
	Cout=> Carry( 	3214	),
	S=> E(	3163	));
			
  U3215	: Soma_AMA3_1 PORT MAP(
	A=> C(	3279	),
	B=>E(	3102	),
	Cin=> Carry( 	3214	),
	Cout=> Carry( 	3215	),
	S=> E(	3164	));
			
  U3216	: Soma_AMA3_1 PORT MAP(
	A=> C(	3280	),
	B=>E(	3103	),
	Cin=> Carry( 	3215	),
	Cout=> Carry( 	3216	),
	S=> E(	3165	));
			
  U3217	: Soma_AMA3_1 PORT MAP(
	A=> C(	3281	),
	B=>E(	3104	),
	Cin=> Carry( 	3216	),
	Cout=> Carry( 	3217	),
	S=> E(	3166	));
			
  U3218	: Soma_AMA3_1 PORT MAP(
	A=> C(	3282	),
	B=>E(	3105	),
	Cin=> Carry( 	3217	),
	Cout=> Carry( 	3218	),
	S=> E(	3167	));
			
  U3219	: Soma_AMA3_1 PORT MAP(
	A=> C(	3283	),
	B=>E(	3106	),
	Cin=> Carry( 	3218	),
	Cout=> Carry( 	3219	),
	S=> E(	3168	));
			
  U3220	: Soma_AMA3_1 PORT MAP(
	A=> C(	3284	),
	B=>E(	3107	),
	Cin=> Carry( 	3219	),
	Cout=> Carry( 	3220	),
	S=> E(	3169	));
			
  U3221	: Soma_AMA3_1 PORT MAP(
	A=> C(	3285	),
	B=>E(	3108	),
	Cin=> Carry( 	3220	),
	Cout=> Carry( 	3221	),
	S=> E(	3170	));
			
  U3222	: Soma_AMA3_1 PORT MAP(
	A=> C(	3286	),
	B=>E(	3109	),
	Cin=> Carry( 	3221	),
	Cout=> Carry( 	3222	),
	S=> E(	3171	));
			
  U3223	: Soma_AMA3_1 PORT MAP(
	A=> C(	3287	),
	B=>E(	3110	),
	Cin=> Carry( 	3222	),
	Cout=> Carry( 	3223	),
	S=> E(	3172	));
			
  U3224	: Soma_AMA3_1 PORT MAP(
	A=> C(	3288	),
	B=>E(	3111	),
	Cin=> Carry( 	3223	),
	Cout=> Carry( 	3224	),
	S=> E(	3173	));
			
  U3225	: Soma_AMA3_1 PORT MAP(
	A=> C(	3289	),
	B=>E(	3112	),
	Cin=> Carry( 	3224	),
	Cout=> Carry( 	3225	),
	S=> E(	3174	));
			
  U3226	: Soma_AMA3_1 PORT MAP(
	A=> C(	3290	),
	B=>E(	3113	),
	Cin=> Carry( 	3225	),
	Cout=> Carry( 	3226	),
	S=> E(	3175	));
			
  U3227	: Soma_AMA3_1 PORT MAP(
	A=> C(	3291	),
	B=>E(	3114	),
	Cin=> Carry( 	3226	),
	Cout=> Carry( 	3227	),
	S=> E(	3176	));
			
  U3228	: Soma_AMA3_1 PORT MAP(
	A=> C(	3292	),
	B=>E(	3115	),
	Cin=> Carry( 	3227	),
	Cout=> Carry( 	3228	),
	S=> E(	3177	));
			
  U3229	: Soma_AMA3_1 PORT MAP(
	A=> C(	3293	),
	B=>E(	3116	),
	Cin=> Carry( 	3228	),
	Cout=> Carry( 	3229	),
	S=> E(	3178	));
			
  U3230	: Soma_AMA3_1 PORT MAP(
	A=> C(	3294	),
	B=>E(	3117	),
	Cin=> Carry( 	3229	),
	Cout=> Carry( 	3230	),
	S=> E(	3179	));
			
  U3231	: Soma_AMA3_1 PORT MAP(
	A=> C(	3295	),
	B=>E(	3118	),
	Cin=> Carry( 	3230	),
	Cout=> Carry( 	3231	),
	S=> E(	3180	));
			
  U3232	: Soma_AMA3_1 PORT MAP(
	A=> C(	3296	),
	B=>E(	3119	),
	Cin=> Carry( 	3231	),
	Cout=> Carry( 	3232	),
	S=> E(	3181	));
			
  U3233	: Soma_AMA3_1 PORT MAP(
	A=> C(	3297	),
	B=>E(	3120	),
	Cin=> Carry( 	3232	),
	Cout=> Carry( 	3233	),
	S=> E(	3182	));
			
  U3234	: Soma_AMA3_1 PORT MAP(
	A=> C(	3298	),
	B=>E(	3121	),
	Cin=> Carry( 	3233	),
	Cout=> Carry( 	3234	),
	S=> E(	3183	));
			
  U3235	: Soma_AMA3_1 PORT MAP(
	A=> C(	3299	),
	B=>E(	3122	),
	Cin=> Carry( 	3234	),
	Cout=> Carry( 	3235	),
	S=> E(	3184	));
			
  U3236	: Soma_AMA3_1 PORT MAP(
	A=> C(	3300	),
	B=>E(	3123	),
	Cin=> Carry( 	3235	),
	Cout=> Carry( 	3236	),
	S=> E(	3185	));
			
  U3237	: Soma_AMA3_1 PORT MAP(
	A=> C(	3301	),
	B=>E(	3124	),
	Cin=> Carry( 	3236	),
	Cout=> Carry( 	3237	),
	S=> E(	3186	));
			
  U3238	: Soma_AMA3_1 PORT MAP(
	A=> C(	3302	),
	B=>E(	3125	),
	Cin=> Carry( 	3237	),
	Cout=> Carry( 	3238	),
	S=> E(	3187	));
			
  U3239	: Soma_AMA3_1 PORT MAP(
	A=> C(	3303	),
	B=>E(	3126	),
	Cin=> Carry( 	3238	),
	Cout=> Carry( 	3239	),
	S=> E(	3188	));
			
  U3240	: Soma_AMA3_1 PORT MAP(
	A=> C(	3304	),
	B=>E(	3127	),
	Cin=> Carry( 	3239	),
	Cout=> Carry( 	3240	),
	S=> E(	3189	));
			
  U3241	: Soma_AMA3_1 PORT MAP(
	A=> C(	3305	),
	B=>E(	3128	),
	Cin=> Carry( 	3240	),
	Cout=> Carry( 	3241	),
	S=> E(	3190	));
			
  U3242	: Soma_AMA3_1 PORT MAP(
	A=> C(	3306	),
	B=>E(	3129	),
	Cin=> Carry( 	3241	),
	Cout=> Carry( 	3242	),
	S=> E(	3191	));
			
  U3243	: Soma_AMA3_1 PORT MAP(
	A=> C(	3307	),
	B=>E(	3130	),
	Cin=> Carry( 	3242	),
	Cout=> Carry( 	3243	),
	S=> E(	3192	));
			
  U3244	: Soma_AMA3_1 PORT MAP(
	A=> C(	3308	),
	B=>E(	3131	),
	Cin=> Carry( 	3243	),
	Cout=> Carry( 	3244	),
	S=> E(	3193	));
			
  U3245	: Soma_AMA3_1 PORT MAP(
	A=> C(	3309	),
	B=>E(	3132	),
	Cin=> Carry( 	3244	),
	Cout=> Carry( 	3245	),
	S=> E(	3194	));
			
  U3246	: Soma_AMA3_1 PORT MAP(
	A=> C(	3310	),
	B=>E(	3133	),
	Cin=> Carry( 	3245	),
	Cout=> Carry( 	3246	),
	S=> E(	3195	));
			
  U3247	: Soma_AMA3_1 PORT MAP(
	A=> C(	3311	),
	B=>E(	3134	),
	Cin=> Carry( 	3246	),
	Cout=> Carry( 	3247	),
	S=> E(	3196	));
			
  U3248	: Soma_AMA3_1 PORT MAP(
	A=> C(	3312	),
	B=>E(	3135	),
	Cin=> Carry( 	3247	),
	Cout=> Carry( 	3248	),
	S=> E(	3197	));
			
  U3249	: Soma_AMA3_1 PORT MAP(
	A=> C(	3313	),
	B=>E(	3136	),
	Cin=> Carry( 	3248	),
	Cout=> Carry( 	3249	),
	S=> E(	3198	));
			
  U3250	: Soma_AMA3_1 PORT MAP(
	A=> C(	3314	),
	B=>E(	3137	),
	Cin=> Carry( 	3249	),
	Cout=> Carry( 	3250	),
	S=> E(	3199	));
			
  U3251	: Soma_AMA3_1 PORT MAP(
	A=> C(	3315	),
	B=>E(	3138	),
	Cin=> Carry( 	3250	),
	Cout=> Carry( 	3251	),
	S=> E(	3200	));
			
  U3252	: Soma_AMA3_1 PORT MAP(
	A=> C(	3316	),
	B=>E(	3139	),
	Cin=> Carry( 	3251	),
	Cout=> Carry( 	3252	),
	S=> E(	3201	));
			
  U3253	: Soma_AMA3_1 PORT MAP(
	A=> C(	3317	),
	B=>E(	3140	),
	Cin=> Carry( 	3252	),
	Cout=> Carry( 	3253	),
	S=> E(	3202	));
			
  U3254	: Soma_AMA3_1 PORT MAP(
	A=> C(	3318	),
	B=>E(	3141	),
	Cin=> Carry( 	3253	),
	Cout=> Carry( 	3254	),
	S=> E(	3203	));
			
  U3255	: Soma_AMA3_1 PORT MAP(
	A=> C(	3319	),
	B=>E(	3142	),
	Cin=> Carry( 	3254	),
	Cout=> Carry( 	3255	),
	S=> E(	3204	));
			
  U3256	: Soma_AMA3_1 PORT MAP(
	A=> C(	3320	),
	B=>E(	3143	),
	Cin=> Carry( 	3255	),
	Cout=> Carry( 	3256	),
	S=> E(	3205	));
			
  U3257	: Soma_AMA3_1 PORT MAP(
	A=> C(	3321	),
	B=>E(	3144	),
	Cin=> Carry( 	3256	),
	Cout=> Carry( 	3257	),
	S=> E(	3206	));
			
  U3258	: Soma_AMA3_1 PORT MAP(
	A=> C(	3322	),
	B=>E(	3145	),
	Cin=> Carry( 	3257	),
	Cout=> Carry( 	3258	),
	S=> E(	3207	));
			
  U3259	: Soma_AMA3_1 PORT MAP(
	A=> C(	3323	),
	B=>E(	3146	),
	Cin=> Carry( 	3258	),
	Cout=> Carry( 	3259	),
	S=> E(	3208	));
			
  U3260	: Soma_AMA3_1 PORT MAP(
	A=> C(	3324	),
	B=>E(	3147	),
	Cin=> Carry( 	3259	),
	Cout=> Carry( 	3260	),
	S=> E(	3209	));
			
  U3261	: Soma_AMA3_1 PORT MAP(
	A=> C(	3325	),
	B=>E(	3148	),
	Cin=> Carry( 	3260	),
	Cout=> Carry( 	3261	),
	S=> E(	3210	));
			
  U3262	: Soma_AMA3_1 PORT MAP(
	A=> C(	3326	),
	B=>E(	3149	),
	Cin=> Carry( 	3261	),
	Cout=> Carry( 	3262	),
	S=> E(	3211	));
			
  U3263	: Soma_AMA3_1 PORT MAP(
	A=> C(	3327	),
	B=>Carry(	3199	),
	Cin=> Carry( 	3262	),
	Cout=> Carry( 	3263	),
	S=> E(	3212	));


			
  U3264	: Soma_AMA3_1 PORT MAP(
	A=> C(	3328	),
	B=>E(	3150	),
	Cin=> '0'	,
	Cout=> Carry( 	3264	),
	S=> R(	52	));
			
  U3265	: Soma_AMA3_1 PORT MAP(
	A=> C(	3329	),
	B=>E(	3151	),
	Cin=> Carry( 	3264	),
	Cout=> Carry( 	3265	),
	S=> E(	3213	));
			
  U3266	: Soma_AMA3_1 PORT MAP(
	A=> C(	3330	),
	B=>E(	3152	),
	Cin=> Carry( 	3265	),
	Cout=> Carry( 	3266	),
	S=> E(	3214	));
			
  U3267	: Soma_AMA3_1 PORT MAP(
	A=> C(	3331	),
	B=>E(	3153	),
	Cin=> Carry( 	3266	),
	Cout=> Carry( 	3267	),
	S=> E(	3215	));
			
  U3268	: Soma_AMA3_1 PORT MAP(
	A=> C(	3332	),
	B=>E(	3154	),
	Cin=> Carry( 	3267	),
	Cout=> Carry( 	3268	),
	S=> E(	3216	));
			
  U3269	: Soma_AMA3_1 PORT MAP(
	A=> C(	3333	),
	B=>E(	3155	),
	Cin=> Carry( 	3268	),
	Cout=> Carry( 	3269	),
	S=> E(	3217	));
			
  U3270	: Soma_AMA3_1 PORT MAP(
	A=> C(	3334	),
	B=>E(	3156	),
	Cin=> Carry( 	3269	),
	Cout=> Carry( 	3270	),
	S=> E(	3218	));
			
  U3271	: Soma_AMA3_1 PORT MAP(
	A=> C(	3335	),
	B=>E(	3157	),
	Cin=> Carry( 	3270	),
	Cout=> Carry( 	3271	),
	S=> E(	3219	));
			
  U3272	: Soma_AMA3_1 PORT MAP(
	A=> C(	3336	),
	B=>E(	3158	),
	Cin=> Carry( 	3271	),
	Cout=> Carry( 	3272	),
	S=> E(	3220	));
			
  U3273	: Soma_AMA3_1 PORT MAP(
	A=> C(	3337	),
	B=>E(	3159	),
	Cin=> Carry( 	3272	),
	Cout=> Carry( 	3273	),
	S=> E(	3221	));
			
  U3274	: Soma_AMA3_1 PORT MAP(
	A=> C(	3338	),
	B=>E(	3160	),
	Cin=> Carry( 	3273	),
	Cout=> Carry( 	3274	),
	S=> E(	3222	));
			
  U3275	: Soma_AMA3_1 PORT MAP(
	A=> C(	3339	),
	B=>E(	3161	),
	Cin=> Carry( 	3274	),
	Cout=> Carry( 	3275	),
	S=> E(	3223	));
			
  U3276	: Soma_AMA3_1 PORT MAP(
	A=> C(	3340	),
	B=>E(	3162	),
	Cin=> Carry( 	3275	),
	Cout=> Carry( 	3276	),
	S=> E(	3224	));
			
  U3277	: Soma_AMA3_1 PORT MAP(
	A=> C(	3341	),
	B=>E(	3163	),
	Cin=> Carry( 	3276	),
	Cout=> Carry( 	3277	),
	S=> E(	3225	));
			
  U3278	: Soma_AMA3_1 PORT MAP(
	A=> C(	3342	),
	B=>E(	3164	),
	Cin=> Carry( 	3277	),
	Cout=> Carry( 	3278	),
	S=> E(	3226	));
			
  U3279	: Soma_AMA3_1 PORT MAP(
	A=> C(	3343	),
	B=>E(	3165	),
	Cin=> Carry( 	3278	),
	Cout=> Carry( 	3279	),
	S=> E(	3227	));
			
  U3280	: Soma_AMA3_1 PORT MAP(
	A=> C(	3344	),
	B=>E(	3166	),
	Cin=> Carry( 	3279	),
	Cout=> Carry( 	3280	),
	S=> E(	3228	));
			
  U3281	: Soma_AMA3_1 PORT MAP(
	A=> C(	3345	),
	B=>E(	3167	),
	Cin=> Carry( 	3280	),
	Cout=> Carry( 	3281	),
	S=> E(	3229	));
			
  U3282	: Soma_AMA3_1 PORT MAP(
	A=> C(	3346	),
	B=>E(	3168	),
	Cin=> Carry( 	3281	),
	Cout=> Carry( 	3282	),
	S=> E(	3230	));
			
  U3283	: Soma_AMA3_1 PORT MAP(
	A=> C(	3347	),
	B=>E(	3169	),
	Cin=> Carry( 	3282	),
	Cout=> Carry( 	3283	),
	S=> E(	3231	));
			
  U3284	: Soma_AMA3_1 PORT MAP(
	A=> C(	3348	),
	B=>E(	3170	),
	Cin=> Carry( 	3283	),
	Cout=> Carry( 	3284	),
	S=> E(	3232	));
			
  U3285	: Soma_AMA3_1 PORT MAP(
	A=> C(	3349	),
	B=>E(	3171	),
	Cin=> Carry( 	3284	),
	Cout=> Carry( 	3285	),
	S=> E(	3233	));
			
  U3286	: Soma_AMA3_1 PORT MAP(
	A=> C(	3350	),
	B=>E(	3172	),
	Cin=> Carry( 	3285	),
	Cout=> Carry( 	3286	),
	S=> E(	3234	));
			
  U3287	: Soma_AMA3_1 PORT MAP(
	A=> C(	3351	),
	B=>E(	3173	),
	Cin=> Carry( 	3286	),
	Cout=> Carry( 	3287	),
	S=> E(	3235	));
			
  U3288	: Soma_AMA3_1 PORT MAP(
	A=> C(	3352	),
	B=>E(	3174	),
	Cin=> Carry( 	3287	),
	Cout=> Carry( 	3288	),
	S=> E(	3236	));
			
  U3289	: Soma_AMA3_1 PORT MAP(
	A=> C(	3353	),
	B=>E(	3175	),
	Cin=> Carry( 	3288	),
	Cout=> Carry( 	3289	),
	S=> E(	3237	));
			
  U3290	: Soma_AMA3_1 PORT MAP(
	A=> C(	3354	),
	B=>E(	3176	),
	Cin=> Carry( 	3289	),
	Cout=> Carry( 	3290	),
	S=> E(	3238	));
			
  U3291	: Soma_AMA3_1 PORT MAP(
	A=> C(	3355	),
	B=>E(	3177	),
	Cin=> Carry( 	3290	),
	Cout=> Carry( 	3291	),
	S=> E(	3239	));
			
  U3292	: Soma_AMA3_1 PORT MAP(
	A=> C(	3356	),
	B=>E(	3178	),
	Cin=> Carry( 	3291	),
	Cout=> Carry( 	3292	),
	S=> E(	3240	));
			
  U3293	: Soma_AMA3_1 PORT MAP(
	A=> C(	3357	),
	B=>E(	3179	),
	Cin=> Carry( 	3292	),
	Cout=> Carry( 	3293	),
	S=> E(	3241	));
			
  U3294	: Soma_AMA3_1 PORT MAP(
	A=> C(	3358	),
	B=>E(	3180	),
	Cin=> Carry( 	3293	),
	Cout=> Carry( 	3294	),
	S=> E(	3242	));
			
  U3295	: Soma_AMA3_1 PORT MAP(
	A=> C(	3359	),
	B=>E(	3181	),
	Cin=> Carry( 	3294	),
	Cout=> Carry( 	3295	),
	S=> E(	3243	));
			
  U3296	: Soma_AMA3_1 PORT MAP(
	A=> C(	3360	),
	B=>E(	3182	),
	Cin=> Carry( 	3295	),
	Cout=> Carry( 	3296	),
	S=> E(	3244	));
			
  U3297	: Soma_AMA3_1 PORT MAP(
	A=> C(	3361	),
	B=>E(	3183	),
	Cin=> Carry( 	3296	),
	Cout=> Carry( 	3297	),
	S=> E(	3245	));
			
  U3298	: Soma_AMA3_1 PORT MAP(
	A=> C(	3362	),
	B=>E(	3184	),
	Cin=> Carry( 	3297	),
	Cout=> Carry( 	3298	),
	S=> E(	3246	));
			
  U3299	: Soma_AMA3_1 PORT MAP(
	A=> C(	3363	),
	B=>E(	3185	),
	Cin=> Carry( 	3298	),
	Cout=> Carry( 	3299	),
	S=> E(	3247	));
			
  U3300	: Soma_AMA3_1 PORT MAP(
	A=> C(	3364	),
	B=>E(	3186	),
	Cin=> Carry( 	3299	),
	Cout=> Carry( 	3300	),
	S=> E(	3248	));
			
  U3301	: Soma_AMA3_1 PORT MAP(
	A=> C(	3365	),
	B=>E(	3187	),
	Cin=> Carry( 	3300	),
	Cout=> Carry( 	3301	),
	S=> E(	3249	));
			
  U3302	: Soma_AMA3_1 PORT MAP(
	A=> C(	3366	),
	B=>E(	3188	),
	Cin=> Carry( 	3301	),
	Cout=> Carry( 	3302	),
	S=> E(	3250	));
			
  U3303	: Soma_AMA3_1 PORT MAP(
	A=> C(	3367	),
	B=>E(	3189	),
	Cin=> Carry( 	3302	),
	Cout=> Carry( 	3303	),
	S=> E(	3251	));
			
  U3304	: Soma_AMA3_1 PORT MAP(
	A=> C(	3368	),
	B=>E(	3190	),
	Cin=> Carry( 	3303	),
	Cout=> Carry( 	3304	),
	S=> E(	3252	));
			
  U3305	: Soma_AMA3_1 PORT MAP(
	A=> C(	3369	),
	B=>E(	3191	),
	Cin=> Carry( 	3304	),
	Cout=> Carry( 	3305	),
	S=> E(	3253	));
			
  U3306	: Soma_AMA3_1 PORT MAP(
	A=> C(	3370	),
	B=>E(	3192	),
	Cin=> Carry( 	3305	),
	Cout=> Carry( 	3306	),
	S=> E(	3254	));
			
  U3307	: Soma_AMA3_1 PORT MAP(
	A=> C(	3371	),
	B=>E(	3193	),
	Cin=> Carry( 	3306	),
	Cout=> Carry( 	3307	),
	S=> E(	3255	));
			
  U3308	: Soma_AMA3_1 PORT MAP(
	A=> C(	3372	),
	B=>E(	3194	),
	Cin=> Carry( 	3307	),
	Cout=> Carry( 	3308	),
	S=> E(	3256	));
			
  U3309	: Soma_AMA3_1 PORT MAP(
	A=> C(	3373	),
	B=>E(	3195	),
	Cin=> Carry( 	3308	),
	Cout=> Carry( 	3309	),
	S=> E(	3257	));
			
  U3310	: Soma_AMA3_1 PORT MAP(
	A=> C(	3374	),
	B=>E(	3196	),
	Cin=> Carry( 	3309	),
	Cout=> Carry( 	3310	),
	S=> E(	3258	));
			
  U3311	: Soma_AMA3_1 PORT MAP(
	A=> C(	3375	),
	B=>E(	3197	),
	Cin=> Carry( 	3310	),
	Cout=> Carry( 	3311	),
	S=> E(	3259	));
			
  U3312	: Soma_AMA3_1 PORT MAP(
	A=> C(	3376	),
	B=>E(	3198	),
	Cin=> Carry( 	3311	),
	Cout=> Carry( 	3312	),
	S=> E(	3260	));
			
  U3313	: Soma_AMA3_1 PORT MAP(
	A=> C(	3377	),
	B=>E(	3199	),
	Cin=> Carry( 	3312	),
	Cout=> Carry( 	3313	),
	S=> E(	3261	));
			
  U3314	: Soma_AMA3_1 PORT MAP(
	A=> C(	3378	),
	B=>E(	3200	),
	Cin=> Carry( 	3313	),
	Cout=> Carry( 	3314	),
	S=> E(	3262	));
			
  U3315	: Soma_AMA3_1 PORT MAP(
	A=> C(	3379	),
	B=>E(	3201	),
	Cin=> Carry( 	3314	),
	Cout=> Carry( 	3315	),
	S=> E(	3263	));
			
  U3316	: Soma_AMA3_1 PORT MAP(
	A=> C(	3380	),
	B=>E(	3202	),
	Cin=> Carry( 	3315	),
	Cout=> Carry( 	3316	),
	S=> E(	3264	));
			
  U3317	: Soma_AMA3_1 PORT MAP(
	A=> C(	3381	),
	B=>E(	3203	),
	Cin=> Carry( 	3316	),
	Cout=> Carry( 	3317	),
	S=> E(	3265	));
			
  U3318	: Soma_AMA3_1 PORT MAP(
	A=> C(	3382	),
	B=>E(	3204	),
	Cin=> Carry( 	3317	),
	Cout=> Carry( 	3318	),
	S=> E(	3266	));
			
  U3319	: Soma_AMA3_1 PORT MAP(
	A=> C(	3383	),
	B=>E(	3205	),
	Cin=> Carry( 	3318	),
	Cout=> Carry( 	3319	),
	S=> E(	3267	));
			
  U3320	: Soma_AMA3_1 PORT MAP(
	A=> C(	3384	),
	B=>E(	3206	),
	Cin=> Carry( 	3319	),
	Cout=> Carry( 	3320	),
	S=> E(	3268	));
			
  U3321	: Soma_AMA3_1 PORT MAP(
	A=> C(	3385	),
	B=>E(	3207	),
	Cin=> Carry( 	3320	),
	Cout=> Carry( 	3321	),
	S=> E(	3269	));
			
  U3322	: Soma_AMA3_1 PORT MAP(
	A=> C(	3386	),
	B=>E(	3208	),
	Cin=> Carry( 	3321	),
	Cout=> Carry( 	3322	),
	S=> E(	3270	));
			
  U3323	: Soma_AMA3_1 PORT MAP(
	A=> C(	3387	),
	B=>E(	3209	),
	Cin=> Carry( 	3322	),
	Cout=> Carry( 	3323	),
	S=> E(	3271	));
			
  U3324	: Soma_AMA3_1 PORT MAP(
	A=> C(	3388	),
	B=>E(	3210	),
	Cin=> Carry( 	3323	),
	Cout=> Carry( 	3324	),
	S=> E(	3272	));
			
  U3325	: Soma_AMA3_1 PORT MAP(
	A=> C(	3389	),
	B=>E(	3211	),
	Cin=> Carry( 	3324	),
	Cout=> Carry( 	3325	),
	S=> E(	3273	));
			
  U3326	: Soma_AMA3_1 PORT MAP(
	A=> C(	3390	),
	B=>E(	3212	),
	Cin=> Carry( 	3325	),
	Cout=> Carry( 	3326	),
	S=> E(	3274	));
			
  U3327	: Soma_AMA3_1 PORT MAP(
	A=> C(	3391	),
	B=>Carry(	3263	),
	Cin=> Carry( 	3326	),
	Cout=> Carry( 	3327	),
	S=> E(	3275	));

			
  U3328	: Soma_AMA3_1 PORT MAP(
	A=> C(	3392	),
	B=>E(	3213	),
	Cin=> '0'	,
	Cout=> Carry( 	3328	),
	S=> R(	53	));
			
  U3329	: Soma_AMA3_1 PORT MAP(
	A=> C(	3393	),
	B=>E(	3214	),
	Cin=> Carry( 	3328	),
	Cout=> Carry( 	3329	),
	S=> E(	3276	));
			
  U3330	: Soma_AMA3_1 PORT MAP(
	A=> C(	3394	),
	B=>E(	3215	),
	Cin=> Carry( 	3329	),
	Cout=> Carry( 	3330	),
	S=> E(	3277	));
			
  U3331	: Soma_AMA3_1 PORT MAP(
	A=> C(	3395	),
	B=>E(	3216	),
	Cin=> Carry( 	3330	),
	Cout=> Carry( 	3331	),
	S=> E(	3278	));
			
  U3332	: Soma_AMA3_1 PORT MAP(
	A=> C(	3396	),
	B=>E(	3217	),
	Cin=> Carry( 	3331	),
	Cout=> Carry( 	3332	),
	S=> E(	3279	));
			
  U3333	: Soma_AMA3_1 PORT MAP(
	A=> C(	3397	),
	B=>E(	3218	),
	Cin=> Carry( 	3332	),
	Cout=> Carry( 	3333	),
	S=> E(	3280	));
			
  U3334	: Soma_AMA3_1 PORT MAP(
	A=> C(	3398	),
	B=>E(	3219	),
	Cin=> Carry( 	3333	),
	Cout=> Carry( 	3334	),
	S=> E(	3281	));
			
  U3335	: Soma_AMA3_1 PORT MAP(
	A=> C(	3399	),
	B=>E(	3220	),
	Cin=> Carry( 	3334	),
	Cout=> Carry( 	3335	),
	S=> E(	3282	));
			
  U3336	: Soma_AMA3_1 PORT MAP(
	A=> C(	3400	),
	B=>E(	3221	),
	Cin=> Carry( 	3335	),
	Cout=> Carry( 	3336	),
	S=> E(	3283	));
			
  U3337	: Soma_AMA3_1 PORT MAP(
	A=> C(	3401	),
	B=>E(	3222	),
	Cin=> Carry( 	3336	),
	Cout=> Carry( 	3337	),
	S=> E(	3284	));
			
  U3338	: Soma_AMA3_1 PORT MAP(
	A=> C(	3402	),
	B=>E(	3223	),
	Cin=> Carry( 	3337	),
	Cout=> Carry( 	3338	),
	S=> E(	3285	));
			
  U3339	: Soma_AMA3_1 PORT MAP(
	A=> C(	3403	),
	B=>E(	3224	),
	Cin=> Carry( 	3338	),
	Cout=> Carry( 	3339	),
	S=> E(	3286	));
			
  U3340	: Soma_AMA3_1 PORT MAP(
	A=> C(	3404	),
	B=>E(	3225	),
	Cin=> Carry( 	3339	),
	Cout=> Carry( 	3340	),
	S=> E(	3287	));
			
  U3341	: Soma_AMA3_1 PORT MAP(
	A=> C(	3405	),
	B=>E(	3226	),
	Cin=> Carry( 	3340	),
	Cout=> Carry( 	3341	),
	S=> E(	3288	));
			
  U3342	: Soma_AMA3_1 PORT MAP(
	A=> C(	3406	),
	B=>E(	3227	),
	Cin=> Carry( 	3341	),
	Cout=> Carry( 	3342	),
	S=> E(	3289	));
			
  U3343	: Soma_AMA3_1 PORT MAP(
	A=> C(	3407	),
	B=>E(	3228	),
	Cin=> Carry( 	3342	),
	Cout=> Carry( 	3343	),
	S=> E(	3290	));
 			
  U3344	: Soma_AMA3_1 PORT MAP(
	A=> C(	3408	),
	B=>E(	3229	),
	Cin=> Carry( 	3343	),
	Cout=> Carry( 	3344	),
	S=> E(	3291	));
			
  U3345	: Soma_AMA3_1 PORT MAP(
	A=> C(	3409	),
	B=>E(	3230	),
	Cin=> Carry( 	3344	),
	Cout=> Carry( 	3345	),
	S=> E(	3292	));
			
  U3346	: Soma_AMA3_1 PORT MAP(
	A=> C(	3410	),
	B=>E(	3231	),
	Cin=> Carry( 	3345	),
	Cout=> Carry( 	3346	),
	S=> E(	3293	));
			
  U3347	: Soma_AMA3_1 PORT MAP(
	A=> C(	3411	),
	B=>E(	3232	),
	Cin=> Carry( 	3346	),
	Cout=> Carry( 	3347	),
	S=> E(	3294	));
			
  U3348	: Soma_AMA3_1 PORT MAP(
	A=> C(	3412	),
	B=>E(	3233	),
	Cin=> Carry( 	3347	),
	Cout=> Carry( 	3348	),
	S=> E(	3295	));
			
  U3349	: Soma_AMA3_1 PORT MAP(
	A=> C(	3413	),
	B=>E(	3234	),
	Cin=> Carry( 	3348	),
	Cout=> Carry( 	3349	),
	S=> E(	3296	));
			
  U3350	: Soma_AMA3_1 PORT MAP(
	A=> C(	3414	),
	B=>E(	3235	),
	Cin=> Carry( 	3349	),
	Cout=> Carry( 	3350	),
	S=> E(	3297	));
			
  U3351	: Soma_AMA3_1 PORT MAP(
	A=> C(	3415	),
	B=>E(	3236	),
	Cin=> Carry( 	3350	),
	Cout=> Carry( 	3351	),
	S=> E(	3298	));
			
  U3352	: Soma_AMA3_1 PORT MAP(
	A=> C(	3416	),
	B=>E(	3237	),
	Cin=> Carry( 	3351	),
	Cout=> Carry( 	3352	),
	S=> E(	3299	));
			
  U3353	: Soma_AMA3_1 PORT MAP(
	A=> C(	3417	),
	B=>E(	3238	),
	Cin=> Carry( 	3352	),
	Cout=> Carry( 	3353	),
	S=> E(	3300	));
			
  U3354	: Soma_AMA3_1 PORT MAP(
	A=> C(	3418	),
	B=>E(	3239	),
	Cin=> Carry( 	3353	),
	Cout=> Carry( 	3354	),
	S=> E(	3301	));
			
  U3355	: Soma_AMA3_1 PORT MAP(
	A=> C(	3419	),
	B=>E(	3240	),
	Cin=> Carry( 	3354	),
	Cout=> Carry( 	3355	),
	S=> E(	3302	));
			
  U3356	: Soma_AMA3_1 PORT MAP(
	A=> C(	3420	),
	B=>E(	3241	),
	Cin=> Carry( 	3355	),
	Cout=> Carry( 	3356	),
	S=> E(	3303	));
			
  U3357	: Soma_AMA3_1 PORT MAP(
	A=> C(	3421	),
	B=>E(	3242	),
	Cin=> Carry( 	3356	),
	Cout=> Carry( 	3357	),
	S=> E(	3304	));
			
  U3358	: Soma_AMA3_1 PORT MAP(
	A=> C(	3422	),
	B=>E(	3243	),
	Cin=> Carry( 	3357	),
	Cout=> Carry( 	3358	),
	S=> E(	3305	));
			
  U3359	: Soma_AMA3_1 PORT MAP(
	A=> C(	3423	),
	B=>E(	3244	),
	Cin=> Carry( 	3358	),
	Cout=> Carry( 	3359	),
	S=> E(	3306	));
			
  U3360	: Soma_AMA3_1 PORT MAP(
	A=> C(	3424	),
	B=>E(	3245	),
	Cin=> Carry( 	3359	),
	Cout=> Carry( 	3360	),
	S=> E(	3307	));
			
  U3361	: Soma_AMA3_1 PORT MAP(
	A=> C(	3425	),
	B=>E(	3246	),
	Cin=> Carry( 	3360	),
	Cout=> Carry( 	3361	),
	S=> E(	3308	));
			
  U3362	: Soma_AMA3_1 PORT MAP(
	A=> C(	3426	),
	B=>E(	3247	),
	Cin=> Carry( 	3361	),
	Cout=> Carry( 	3362	),
	S=> E(	3309	));
			
  U3363	: Soma_AMA3_1 PORT MAP(
	A=> C(	3427	),
	B=>E(	3248	),
	Cin=> Carry( 	3362	),
	Cout=> Carry( 	3363	),
	S=> E(	3310	));
			
  U3364	: Soma_AMA3_1 PORT MAP(
	A=> C(	3428	),
	B=>E(	3249	),
	Cin=> Carry( 	3363	),
	Cout=> Carry( 	3364	),
	S=> E(	3311	));
			
  U3365	: Soma_AMA3_1 PORT MAP(
	A=> C(	3429	),
	B=>E(	3250	),
	Cin=> Carry( 	3364	),
	Cout=> Carry( 	3365	),
	S=> E(	3312	));
			
  U3366	: Soma_AMA3_1 PORT MAP(
	A=> C(	3430	),
	B=>E(	3251	),
	Cin=> Carry( 	3365	),
	Cout=> Carry( 	3366	),
	S=> E(	3313	));
			
  U3367	: Soma_AMA3_1 PORT MAP(
	A=> C(	3431	),
	B=>E(	3252	),
	Cin=> Carry( 	3366	),
	Cout=> Carry( 	3367	),
	S=> E(	3314	));
			
  U3368	: Soma_AMA3_1 PORT MAP(
	A=> C(	3432	),
	B=>E(	3253	),
	Cin=> Carry( 	3367	),
	Cout=> Carry( 	3368	),
	S=> E(	3315	));
			
  U3369	: Soma_AMA3_1 PORT MAP(
	A=> C(	3433	),
	B=>E(	3254	),
	Cin=> Carry( 	3368	),
	Cout=> Carry( 	3369	),
	S=> E(	3316	));
			
  U3370	: Soma_AMA3_1 PORT MAP(
	A=> C(	3434	),
	B=>E(	3255	),
	Cin=> Carry( 	3369	),
	Cout=> Carry( 	3370	),
	S=> E(	3317	));
			
  U3371	: Soma_AMA3_1 PORT MAP(
	A=> C(	3435	),
	B=>E(	3256	),
	Cin=> Carry( 	3370	),
	Cout=> Carry( 	3371	),
	S=> E(	3318	));
			
  U3372	: Soma_AMA3_1 PORT MAP(
	A=> C(	3436	),
	B=>E(	3257	),
	Cin=> Carry( 	3371	),
	Cout=> Carry( 	3372	),
	S=> E(	3319	));
			
  U3373	: Soma_AMA3_1 PORT MAP(
	A=> C(	3437	),
	B=>E(	3258	),
	Cin=> Carry( 	3372	),
	Cout=> Carry( 	3373	),
	S=> E(	3320	));
			
  U3374	: Soma_AMA3_1 PORT MAP(
	A=> C(	3438	),
	B=>E(	3259	),
	Cin=> Carry( 	3373	),
	Cout=> Carry( 	3374	),
	S=> E(	3321	));
			
  U3375	: Soma_AMA3_1 PORT MAP(
	A=> C(	3439	),
	B=>E(	3260	),
	Cin=> Carry( 	3374	),
	Cout=> Carry( 	3375	),
	S=> E(	3322	));
			
  U3376	: Soma_AMA3_1 PORT MAP(
	A=> C(	3440	),
	B=>E(	3261	),
	Cin=> Carry( 	3375	),
	Cout=> Carry( 	3376	),
	S=> E(	3323	));
			
  U3377	: Soma_AMA3_1 PORT MAP(
	A=> C(	3441	),
	B=>E(	3262	),
	Cin=> Carry( 	3376	),
	Cout=> Carry( 	3377	),
	S=> E(	3324	));
			
  U3378	: Soma_AMA3_1 PORT MAP(
	A=> C(	3442	),
	B=>E(	3263	),
	Cin=> Carry( 	3377	),
	Cout=> Carry( 	3378	),
	S=> E(	3325	));
			
  U3379	: Soma_AMA3_1 PORT MAP(
	A=> C(	3443	),
	B=>E(	3264	),
	Cin=> Carry( 	3378	),
	Cout=> Carry( 	3379	),
	S=> E(	3326	));
			
  U3380	: Soma_AMA3_1 PORT MAP(
	A=> C(	3444	),
	B=>E(	3265	),
	Cin=> Carry( 	3379	),
	Cout=> Carry( 	3380	),
	S=> E(	3327	));
			
  U3381	: Soma_AMA3_1 PORT MAP(
	A=> C(	3445	),
	B=>E(	3266	),
	Cin=> Carry( 	3380	),
	Cout=> Carry( 	3381	),
	S=> E(	3328	));
			
  U3382	: Soma_AMA3_1 PORT MAP(
	A=> C(	3446	),
	B=>E(	3267	),
	Cin=> Carry( 	3381	),
	Cout=> Carry( 	3382	),
	S=> E(	3329	));
			
  U3383	: Soma_AMA3_1 PORT MAP(
	A=> C(	3447	),
	B=>E(	3268	),
	Cin=> Carry( 	3382	),
	Cout=> Carry( 	3383	),
	S=> E(	3330	));
			
  U3384	: Soma_AMA3_1 PORT MAP(
	A=> C(	3448	),
	B=>E(	3269	),
	Cin=> Carry( 	3383	),
	Cout=> Carry( 	3384	),
	S=> E(	3331	));
			
  U3385	: Soma_AMA3_1 PORT MAP(
	A=> C(	3449	),
	B=>E(	3270	),
	Cin=> Carry( 	3384	),
	Cout=> Carry( 	3385	),
	S=> E(	3332	));
			
  U3386	: Soma_AMA3_1 PORT MAP(
	A=> C(	3450	),
	B=>E(	3271	),
	Cin=> Carry( 	3385	),
	Cout=> Carry( 	3386	),
	S=> E(	3333	));
			
  U3387	: Soma_AMA3_1 PORT MAP(
	A=> C(	3451	),
	B=>E(	3272	),
	Cin=> Carry( 	3386	),
	Cout=> Carry( 	3387	),
	S=> E(	3334	));
			
  U3388	: Soma_AMA3_1 PORT MAP(
	A=> C(	3452	),
	B=>E(	3273	),
	Cin=> Carry( 	3387	),
	Cout=> Carry( 	3388	),
	S=> E(	3335	));
			
  U3389	: Soma_AMA3_1 PORT MAP(
	A=> C(	3453	),
	B=>E(	3274	),
	Cin=> Carry( 	3388	),
	Cout=> Carry( 	3389	),
	S=> E(	3336	));
			
  U3390	: Soma_AMA3_1 PORT MAP(
	A=> C(	3454	),
	B=>E(	3275	),
	Cin=> Carry( 	3389	),
	Cout=> Carry( 	3390	),
	S=> E(	3337	));
			
  U3391	: Soma_AMA3_1 PORT MAP(
	A=> C(	3455	),
	B=>Carry(	3327	),
	Cin=> Carry( 	3390	),
	Cout=> Carry( 	3391	),
	S=> E(	3338	));
			
  U3392	: Soma_AMA3_1 PORT MAP(
	A=> C(	3456	),
	B=>E(	3276	),
	Cin=> '0'	,
	Cout=> Carry( 	3392	),
	S=> R(	54	));
			
  U3393	: Soma_AMA3_1 PORT MAP(
	A=> C(	3457	),
	B=>E(	3277	),
	Cin=> Carry( 	3392	),
	Cout=> Carry( 	3393	),
	S=> E(	3339	));
			
  U3394	: Soma_AMA3_1 PORT MAP(
	A=> C(	3458	),
	B=>E(	3278	),
	Cin=> Carry( 	3393	),
	Cout=> Carry( 	3394	),
	S=> E(	3340	));
			
  U3395	: Soma_AMA3_1 PORT MAP(
	A=> C(	3459	),
	B=>E(	3279	),
	Cin=> Carry( 	3394	),
	Cout=> Carry( 	3395	),
	S=> E(	3341	));
			
  U3396	: Soma_AMA3_1 PORT MAP(
	A=> C(	3460	),
	B=>E(	3280	),
	Cin=> Carry( 	3395	),
	Cout=> Carry( 	3396	),
	S=> E(	3342	));
			
  U3397	: Soma_AMA3_1 PORT MAP(
	A=> C(	3461	),
	B=>E(	3281	),
	Cin=> Carry( 	3396	),
	Cout=> Carry( 	3397	),
	S=> E(	3343	));
			
  U3398	: Soma_AMA3_1 PORT MAP(
	A=> C(	3462	),
	B=>E(	3282	),
	Cin=> Carry( 	3397	),
	Cout=> Carry( 	3398	),
	S=> E(	3344	));
			
  U3399	: Soma_AMA3_1 PORT MAP(
	A=> C(	3463	),
	B=>E(	3283	),
	Cin=> Carry( 	3398	),
	Cout=> Carry( 	3399	),
	S=> E(	3345	));
			
  U3400	: Soma_AMA3_1 PORT MAP(
	A=> C(	3464	),
	B=>E(	3284	),
	Cin=> Carry( 	3399	),
	Cout=> Carry( 	3400	),
	S=> E(	3346	));
			
  U3401	: Soma_AMA3_1 PORT MAP(
	A=> C(	3465	),
	B=>E(	3285	),
	Cin=> Carry( 	3400	),
	Cout=> Carry( 	3401	),
	S=> E(	3347	));
			
  U3402	: Soma_AMA3_1 PORT MAP(
	A=> C(	3466	),
	B=>E(	3286	),
	Cin=> Carry( 	3401	),
	Cout=> Carry( 	3402	),
	S=> E(	3348	));
			
  U3403	: Soma_AMA3_1 PORT MAP(
	A=> C(	3467	),
	B=>E(	3287	),
	Cin=> Carry( 	3402	),
	Cout=> Carry( 	3403	),
	S=> E(	3349	));
			
  U3404	: Soma_AMA3_1 PORT MAP(
	A=> C(	3468	),
	B=>E(	3288	),
	Cin=> Carry( 	3403	),
	Cout=> Carry( 	3404	),
	S=> E(	3350	));
			
  U3405	: Soma_AMA3_1 PORT MAP(
	A=> C(	3469	),
	B=>E(	3289	),
	Cin=> Carry( 	3404	),
	Cout=> Carry( 	3405	),
	S=> E(	3351	));
			
  U3406	: Soma_AMA3_1 PORT MAP(
	A=> C(	3470	),
	B=>E(	3290	),
	Cin=> Carry( 	3405	),
	Cout=> Carry( 	3406	),
	S=> E(	3352	));
			
  U3407	: Soma_AMA3_1 PORT MAP(
	A=> C(	3471	),
	B=>E(	3291	),
	Cin=> Carry( 	3406	),
	Cout=> Carry( 	3407	),
	S=> E(	3353	));
			
  U3408	: Soma_AMA3_1 PORT MAP(
	A=> C(	3472	),
	B=>E(	3292	),
	Cin=> Carry( 	3407	),
	Cout=> Carry( 	3408	),
	S=> E(	3354	));
			
  U3409	: Soma_AMA3_1 PORT MAP(
	A=> C(	3473	),
	B=>E(	3293	),
	Cin=> Carry( 	3408	),
	Cout=> Carry( 	3409	),
	S=> E(	3355	));
			
  U3410	: Soma_AMA3_1 PORT MAP(
	A=> C(	3474	),
	B=>E(	3294	),
	Cin=> Carry( 	3409	),
	Cout=> Carry( 	3410	),
	S=> E(	3356	));
			
  U3411	: Soma_AMA3_1 PORT MAP(
	A=> C(	3475	),
	B=>E(	3295	),
	Cin=> Carry( 	3410	),
	Cout=> Carry( 	3411	),
	S=> E(	3357	));
			
  U3412	: Soma_AMA3_1 PORT MAP(
	A=> C(	3476	),
	B=>E(	3296	),
	Cin=> Carry( 	3411	),
	Cout=> Carry( 	3412	),
	S=> E(	3358	));
			
  U3413	: Soma_AMA3_1 PORT MAP(
	A=> C(	3477	),
	B=>E(	3297	),
	Cin=> Carry( 	3412	),
	Cout=> Carry( 	3413	),
	S=> E(	3359	));
			
  U3414	: Soma_AMA3_1 PORT MAP(
	A=> C(	3478	),
	B=>E(	3298	),
	Cin=> Carry( 	3413	),
	Cout=> Carry( 	3414	),
	S=> E(	3360	));
			
  U3415	: Soma_AMA3_1 PORT MAP(
	A=> C(	3479	),
	B=>E(	3299	),
	Cin=> Carry( 	3414	),
	Cout=> Carry( 	3415	),
	S=> E(	3361	));
			
  U3416	: Soma_AMA3_1 PORT MAP(
	A=> C(	3480	),
	B=>E(	3300	),
	Cin=> Carry( 	3415	),
	Cout=> Carry( 	3416	),
	S=> E(	3362	));
			
  U3417	: Soma_AMA3_1 PORT MAP(
	A=> C(	3481	),
	B=>E(	3301	),
	Cin=> Carry( 	3416	),
	Cout=> Carry( 	3417	),
	S=> E(	3363	));
			
  U3418	: Soma_AMA3_1 PORT MAP(
	A=> C(	3482	),
	B=>E(	3302	),
	Cin=> Carry( 	3417	),
	Cout=> Carry( 	3418	),
	S=> E(	3364	));
			
  U3419	: Soma_AMA3_1 PORT MAP(
	A=> C(	3483	),
	B=>E(	3303	),
	Cin=> Carry( 	3418	),
	Cout=> Carry( 	3419	),
	S=> E(	3365	));
			
  U3420	: Soma_AMA3_1 PORT MAP(
	A=> C(	3484	),
	B=>E(	3304	),
	Cin=> Carry( 	3419	),
	Cout=> Carry( 	3420	),
	S=> E(	3366	));
			
  U3421	: Soma_AMA3_1 PORT MAP(
	A=> C(	3485	),
	B=>E(	3305	),
	Cin=> Carry( 	3420	),
	Cout=> Carry( 	3421	),
	S=> E(	3367	));
			
  U3422	: Soma_AMA3_1 PORT MAP(
	A=> C(	3486	),
	B=>E(	3306	),
	Cin=> Carry( 	3421	),
	Cout=> Carry( 	3422	),
	S=> E(	3368	));
			
  U3423	: Soma_AMA3_1 PORT MAP(
	A=> C(	3487	),
	B=>E(	3307	),
	Cin=> Carry( 	3422	),
	Cout=> Carry( 	3423	),
	S=> E(	3369	));
			
  U3424	: Soma_AMA3_1 PORT MAP(
	A=> C(	3488	),
	B=>E(	3308	),
	Cin=> Carry( 	3423	),
	Cout=> Carry( 	3424	),
	S=> E(	3370	));
			
  U3425	: Soma_AMA3_1 PORT MAP(
	A=> C(	3489	),
	B=>E(	3309	),
	Cin=> Carry( 	3424	),
	Cout=> Carry( 	3425	),
	S=> E(	3371	));
			
  U3426	: Soma_AMA3_1 PORT MAP(
	A=> C(	3490	),
	B=>E(	3310	),
	Cin=> Carry( 	3425	),
	Cout=> Carry( 	3426	),
	S=> E(	3372	));
			
  U3427	: Soma_AMA3_1 PORT MAP(
	A=> C(	3491	),
	B=>E(	3311	),
	Cin=> Carry( 	3426	),
	Cout=> Carry( 	3427	),
	S=> E(	3373	));
			
  U3428	: Soma_AMA3_1 PORT MAP(
	A=> C(	3492	),
	B=>E(	3312	),
	Cin=> Carry( 	3427	),
	Cout=> Carry( 	3428	),
	S=> E(	3374	));
			
  U3429	: Soma_AMA3_1 PORT MAP(
	A=> C(	3493	),
	B=>E(	3313	),
	Cin=> Carry( 	3428	),
	Cout=> Carry( 	3429	),
	S=> E(	3375	));
			
  U3430	: Soma_AMA3_1 PORT MAP(
	A=> C(	3494	),
	B=>E(	3314	),
	Cin=> Carry( 	3429	),
	Cout=> Carry( 	3430	),
	S=> E(	3376	));
			
  U3431	: Soma_AMA3_1 PORT MAP(
	A=> C(	3495	),
	B=>E(	3315	),
	Cin=> Carry( 	3430	),
	Cout=> Carry( 	3431	),
	S=> E(	3377	));
			
  U3432	: Soma_AMA3_1 PORT MAP(
	A=> C(	3496	),
	B=>E(	3316	),
	Cin=> Carry( 	3431	),
	Cout=> Carry( 	3432	),
	S=> E(	3378	));
			
  U3433	: Soma_AMA3_1 PORT MAP(
	A=> C(	3497	),
	B=>E(	3317	),
	Cin=> Carry( 	3432	),
	Cout=> Carry( 	3433	),
	S=> E(	3379	));
			
  U3434	: Soma_AMA3_1 PORT MAP(
	A=> C(	3498	),
	B=>E(	3318	),
	Cin=> Carry( 	3433	),
	Cout=> Carry( 	3434	),
	S=> E(	3380	));
			
  U3435	: Soma_AMA3_1 PORT MAP(
	A=> C(	3499	),
	B=>E(	3319	),
	Cin=> Carry( 	3434	),
	Cout=> Carry( 	3435	),
	S=> E(	3381	));
			
  U3436	: Soma_AMA3_1 PORT MAP(
	A=> C(	3500	),
	B=>E(	3320	),
	Cin=> Carry( 	3435	),
	Cout=> Carry( 	3436	),
	S=> E(	3382	));
			
  U3437	: Soma_AMA3_1 PORT MAP(
	A=> C(	3501	),
	B=>E(	3321	),
	Cin=> Carry( 	3436	),
	Cout=> Carry( 	3437	),
	S=> E(	3383	));
			
  U3438	: Soma_AMA3_1 PORT MAP(
	A=> C(	3502	),
	B=>E(	3322	),
	Cin=> Carry( 	3437	),
	Cout=> Carry( 	3438	),
	S=> E(	3384	));
			
  U3439	: Soma_AMA3_1 PORT MAP(
	A=> C(	3503	),
	B=>E(	3323	),
	Cin=> Carry( 	3438	),
	Cout=> Carry( 	3439	),
	S=> E(	3385	));
			
  U3440	: Soma_AMA3_1 PORT MAP(
	A=> C(	3504	),
	B=>E(	3324	),
	Cin=> Carry( 	3439	),
	Cout=> Carry( 	3440	),
	S=> E(	3386	));
			
  U3441	: Soma_AMA3_1 PORT MAP(
	A=> C(	3505	),
	B=>E(	3325	),
	Cin=> Carry( 	3440	),
	Cout=> Carry( 	3441	),
	S=> E(	3387	));
			
  U3442	: Soma_AMA3_1 PORT MAP(
	A=> C(	3506	),
	B=>E(	3326	),
	Cin=> Carry( 	3441	),
	Cout=> Carry( 	3442	),
	S=> E(	3388	));
			
  U3443	: Soma_AMA3_1 PORT MAP(
	A=> C(	3507	),
	B=>E(	3327	),
	Cin=> Carry( 	3442	),
	Cout=> Carry( 	3443	),
	S=> E(	3389	));
			
  U3444	: Soma_AMA3_1 PORT MAP(
	A=> C(	3508	),
	B=>E(	3328	),
	Cin=> Carry( 	3443	),
	Cout=> Carry( 	3444	),
	S=> E(	3390	));
			
  U3445	: Soma_AMA3_1 PORT MAP(
	A=> C(	3509	),
	B=>E(	3329	),
	Cin=> Carry( 	3444	),
	Cout=> Carry( 	3445	),
	S=> E(	3391	));
			
  U3446	: Soma_AMA3_1 PORT MAP(
	A=> C(	3510	),
	B=>E(	3330	),
	Cin=> Carry( 	3445	),
	Cout=> Carry( 	3446	),
	S=> E(	3392	));
			
  U3447	: Soma_AMA3_1 PORT MAP(
	A=> C(	3511	),
	B=>E(	3331	),
	Cin=> Carry( 	3446	),
	Cout=> Carry( 	3447	),
	S=> E(	3393	));
			
  U3448	: Soma_AMA3_1 PORT MAP(
	A=> C(	3512	),
	B=>E(	3332	),
	Cin=> Carry( 	3447	),
	Cout=> Carry( 	3448	),
	S=> E(	3394	));
			
  U3449	: Soma_AMA3_1 PORT MAP(
	A=> C(	3513	),
	B=>E(	3333	),
	Cin=> Carry( 	3448	),
	Cout=> Carry( 	3449	),
	S=> E(	3395	));
			
  U3450	: Soma_AMA3_1 PORT MAP(
	A=> C(	3514	),
	B=>E(	3334	),
	Cin=> Carry( 	3449	),
	Cout=> Carry( 	3450	),
	S=> E(	3396	));
			
  U3451	: Soma_AMA3_1 PORT MAP(
	A=> C(	3515	),
	B=>E(	3335	),
	Cin=> Carry( 	3450	),
	Cout=> Carry( 	3451	),
	S=> E(	3397	));
			
  U3452	: Soma_AMA3_1 PORT MAP(
	A=> C(	3516	),
	B=>E(	3336	),
	Cin=> Carry( 	3451	),
	Cout=> Carry( 	3452	),
	S=> E(	3398	));
			
  U3453	: Soma_AMA3_1 PORT MAP(
	A=> C(	3517	),
	B=>E(	3337	),
	Cin=> Carry( 	3452	),
	Cout=> Carry( 	3453	),
	S=> E(	3399	));
			
  U3454	: Soma_AMA3_1 PORT MAP(
	A=> C(	3518	),
	B=>E(	3338	),
	Cin=> Carry( 	3453	),
	Cout=> Carry( 	3454	),
	S=> E(	3400	));
			
  U3455	: Soma_AMA3_1 PORT MAP(
	A=> C(	3519	),
	B=>Carry(	3391	),
	Cin=> Carry( 	3454	),
	Cout=> Carry( 	3455	),
	S=> E(	3401	));

			
  U3456	: Soma_AMA3_1 PORT MAP(
	A=> C(	3520	),
	B=>E(	3339	),
	Cin=> '0'	,
	Cout=> Carry( 	3456	),
	S=> R(	55	));
			
  U3457	: Soma_AMA3_1 PORT MAP(
	A=> C(	3521	),
	B=>E(	3340	),
	Cin=> Carry( 	3456	),
	Cout=> Carry( 	3457	),
	S=> E(	3402	));
			
  U3458	: Soma_AMA3_1 PORT MAP(
	A=> C(	3522	),
	B=>E(	3341	),
	Cin=> Carry( 	3457	),
	Cout=> Carry( 	3458	),
	S=> E(	3403	));
			
  U3459	: Soma_AMA3_1 PORT MAP(
	A=> C(	3523	),
	B=>E(	3342	),
	Cin=> Carry( 	3458	),
	Cout=> Carry( 	3459	),
	S=> E(	3404	));
			
  U3460	: Soma_AMA3_1 PORT MAP(
	A=> C(	3524	),
	B=>E(	3343	),
	Cin=> Carry( 	3459	),
	Cout=> Carry( 	3460	),
	S=> E(	3405	));
			
  U3461	: Soma_AMA3_1 PORT MAP(
	A=> C(	3525	),
	B=>E(	3344	),
	Cin=> Carry( 	3460	),
	Cout=> Carry( 	3461	),
	S=> E(	3406	));
			
  U3462	: Soma_AMA3_1 PORT MAP(
	A=> C(	3526	),
	B=>E(	3345	),
	Cin=> Carry( 	3461	),
	Cout=> Carry( 	3462	),
	S=> E(	3407	));
			
  U3463	: Soma_AMA3_1 PORT MAP(
	A=> C(	3527	),
	B=>E(	3346	),
	Cin=> Carry( 	3462	),
	Cout=> Carry( 	3463	),
	S=> E(	3408	));
			
  U3464	: Soma_AMA3_1 PORT MAP(
	A=> C(	3528	),
	B=>E(	3347	),
	Cin=> Carry( 	3463	),
	Cout=> Carry( 	3464	),
	S=> E(	3409	));
			
  U3465	: Soma_AMA3_1 PORT MAP(
	A=> C(	3529	),
	B=>E(	3348	),
	Cin=> Carry( 	3464	),
	Cout=> Carry( 	3465	),
	S=> E(	3410	));
			
  U3466	: Soma_AMA3_1 PORT MAP(
	A=> C(	3530	),
	B=>E(	3349	),
	Cin=> Carry( 	3465	),
	Cout=> Carry( 	3466	),
	S=> E(	3411	));
			
  U3467	: Soma_AMA3_1 PORT MAP(
	A=> C(	3531	),
	B=>E(	3350	),
	Cin=> Carry( 	3466	),
	Cout=> Carry( 	3467	),
	S=> E(	3412	));
			
  U3468	: Soma_AMA3_1 PORT MAP(
	A=> C(	3532	),
	B=>E(	3351	),
	Cin=> Carry( 	3467	),
	Cout=> Carry( 	3468	),
	S=> E(	3413	));
			
  U3469	: Soma_AMA3_1 PORT MAP(
	A=> C(	3533	),
	B=>E(	3352	),
	Cin=> Carry( 	3468	),
	Cout=> Carry( 	3469	),
	S=> E(	3414	));
			
  U3470	: Soma_AMA3_1 PORT MAP(
	A=> C(	3534	),
	B=>E(	3353	),
	Cin=> Carry( 	3469	),
	Cout=> Carry( 	3470	),
	S=> E(	3415	));
			
  U3471	: Soma_AMA3_1 PORT MAP(
	A=> C(	3535	),
	B=>E(	3354	),
	Cin=> Carry( 	3470	),
	Cout=> Carry( 	3471	),
	S=> E(	3416	));
			
  U3472	: Soma_AMA3_1 PORT MAP(
	A=> C(	3536	),
	B=>E(	3355	),
	Cin=> Carry( 	3471	),
	Cout=> Carry( 	3472	),
	S=> E(	3417	));
			
  U3473	: Soma_AMA3_1 PORT MAP(
	A=> C(	3537	),
	B=>E(	3356	),
	Cin=> Carry( 	3472	),
	Cout=> Carry( 	3473	),
	S=> E(	3418	));
			
  U3474	: Soma_AMA3_1 PORT MAP(
	A=> C(	3538	),
	B=>E(	3357	),
	Cin=> Carry( 	3473	),
	Cout=> Carry( 	3474	),
	S=> E(	3419	));
			
  U3475	: Soma_AMA3_1 PORT MAP(
	A=> C(	3539	),
	B=>E(	3358	),
	Cin=> Carry( 	3474	),
	Cout=> Carry( 	3475	),
	S=> E(	3420	));
			
  U3476	: Soma_AMA3_1 PORT MAP(
	A=> C(	3540	),
	B=>E(	3359	),
	Cin=> Carry( 	3475	),
	Cout=> Carry( 	3476	),
	S=> E(	3421	));
			
  U3477	: Soma_AMA3_1 PORT MAP(
	A=> C(	3541	),
	B=>E(	3360	),
	Cin=> Carry( 	3476	),
	Cout=> Carry( 	3477	),
	S=> E(	3422	));
			
  U3478	: Soma_AMA3_1 PORT MAP(
	A=> C(	3542	),
	B=>E(	3361	),
	Cin=> Carry( 	3477	),
	Cout=> Carry( 	3478	),
	S=> E(	3423	));
			
  U3479	: Soma_AMA3_1 PORT MAP(
	A=> C(	3543	),
	B=>E(	3362	),
	Cin=> Carry( 	3478	),
	Cout=> Carry( 	3479	),
	S=> E(	3424	));
			
  U3480	: Soma_AMA3_1 PORT MAP(
	A=> C(	3544	),
	B=>E(	3363	),
	Cin=> Carry( 	3479	),
	Cout=> Carry( 	3480	),
	S=> E(	3425	));
			
  U3481	: Soma_AMA3_1 PORT MAP(
	A=> C(	3545	),
	B=>E(	3364	),
	Cin=> Carry( 	3480	),
	Cout=> Carry( 	3481	),
	S=> E(	3426	));
			
  U3482	: Soma_AMA3_1 PORT MAP(
	A=> C(	3546	),
	B=>E(	3365	),
	Cin=> Carry( 	3481	),
	Cout=> Carry( 	3482	),
	S=> E(	3427	));
			
  U3483	: Soma_AMA3_1 PORT MAP(
	A=> C(	3547	),
	B=>E(	3366	),
	Cin=> Carry( 	3482	),
	Cout=> Carry( 	3483	),
	S=> E(	3428	));
			
  U3484	: Soma_AMA3_1 PORT MAP(
	A=> C(	3548	),
	B=>E(	3367	),
	Cin=> Carry( 	3483	),
	Cout=> Carry( 	3484	),
	S=> E(	3429	));
			
  U3485	: Soma_AMA3_1 PORT MAP(
	A=> C(	3549	),
	B=>E(	3368	),
	Cin=> Carry( 	3484	),
	Cout=> Carry( 	3485	),
	S=> E(	3430	));
			
  U3486	: Soma_AMA3_1 PORT MAP(
	A=> C(	3550	),
	B=>E(	3369	),
	Cin=> Carry( 	3485	),
	Cout=> Carry( 	3486	),
	S=> E(	3431	));
			
  U3487	: Soma_AMA3_1 PORT MAP(
	A=> C(	3551	),
	B=>E(	3370	),
	Cin=> Carry( 	3486	),
	Cout=> Carry( 	3487	),
	S=> E(	3432	));
			
  U3488	: Soma_AMA3_1 PORT MAP(
	A=> C(	3552	),
	B=>E(	3371	),
	Cin=> Carry( 	3487	),
	Cout=> Carry( 	3488	),
	S=> E(	3433	));
			
  U3489	: Soma_AMA3_1 PORT MAP(
	A=> C(	3553	),
	B=>E(	3372	),
	Cin=> Carry( 	3488	),
	Cout=> Carry( 	3489	),
	S=> E(	3434	));
			
  U3490	: Soma_AMA3_1 PORT MAP(
	A=> C(	3554	),
	B=>E(	3373	),
	Cin=> Carry( 	3489	),
	Cout=> Carry( 	3490	),
	S=> E(	3435	));
			
  U3491	: Soma_AMA3_1 PORT MAP(
	A=> C(	3555	),
	B=>E(	3374	),
	Cin=> Carry( 	3490	),
	Cout=> Carry( 	3491	),
	S=> E(	3436	));
			
  U3492	: Soma_AMA3_1 PORT MAP(
	A=> C(	3556	),
	B=>E(	3375	),
	Cin=> Carry( 	3491	),
	Cout=> Carry( 	3492	),
	S=> E(	3437	));
			
  U3493	: Soma_AMA3_1 PORT MAP(
	A=> C(	3557	),
	B=>E(	3376	),
	Cin=> Carry( 	3492	),
	Cout=> Carry( 	3493	),
	S=> E(	3438	));
			
  U3494	: Soma_AMA3_1 PORT MAP(
	A=> C(	3558	),
	B=>E(	3377	),
	Cin=> Carry( 	3493	),
	Cout=> Carry( 	3494	),
	S=> E(	3439	));
			
  U3495	: Soma_AMA3_1 PORT MAP(
	A=> C(	3559	),
	B=>E(	3378	),
	Cin=> Carry( 	3494	),
	Cout=> Carry( 	3495	),
	S=> E(	3440	));
			
  U3496	: Soma_AMA3_1 PORT MAP(
	A=> C(	3560	),
	B=>E(	3379	),
	Cin=> Carry( 	3495	),
	Cout=> Carry( 	3496	),
	S=> E(	3441	));
			
  U3497	: Soma_AMA3_1 PORT MAP(
	A=> C(	3561	),
	B=>E(	3380	),
	Cin=> Carry( 	3496	),
	Cout=> Carry( 	3497	),
	S=> E(	3442	));
			
  U3498	: Soma_AMA3_1 PORT MAP(
	A=> C(	3562	),
	B=>E(	3381	),
	Cin=> Carry( 	3497	),
	Cout=> Carry( 	3498	),
	S=> E(	3443	));
			
  U3499	: Soma_AMA3_1 PORT MAP(
	A=> C(	3563	),
	B=>E(	3382	),
	Cin=> Carry( 	3498	),
	Cout=> Carry( 	3499	),
	S=> E(	3444	));
			
  U3500	: Soma_AMA3_1 PORT MAP(
	A=> C(	3564	),
	B=>E(	3383	),
	Cin=> Carry( 	3499	),
	Cout=> Carry( 	3500	),
	S=> E(	3445	));
			
  U3501	: Soma_AMA3_1 PORT MAP(
	A=> C(	3565	),
	B=>E(	3384	),
	Cin=> Carry( 	3500	),
	Cout=> Carry( 	3501	),
	S=> E(	3446	));
			
  U3502	: Soma_AMA3_1 PORT MAP(
	A=> C(	3566	),
	B=>E(	3385	),
	Cin=> Carry( 	3501	),
	Cout=> Carry( 	3502	),
	S=> E(	3447	));
			
  U3503	: Soma_AMA3_1 PORT MAP(
	A=> C(	3567	),
	B=>E(	3386	),
	Cin=> Carry( 	3502	),
	Cout=> Carry( 	3503	),
	S=> E(	3448	));
			
  U3504	: Soma_AMA3_1 PORT MAP(
	A=> C(	3568	),
	B=>E(	3387	),
	Cin=> Carry( 	3503	),
	Cout=> Carry( 	3504	),
	S=> E(	3449	));
			
  U3505	: Soma_AMA3_1 PORT MAP(
	A=> C(	3569	),
	B=>E(	3388	),
	Cin=> Carry( 	3504	),
	Cout=> Carry( 	3505	),
	S=> E(	3450	));
			
  U3506	: Soma_AMA3_1 PORT MAP(
	A=> C(	3570	),
	B=>E(	3389	),
	Cin=> Carry( 	3505	),
	Cout=> Carry( 	3506	),
	S=> E(	3451	));
			
  U3507	: Soma_AMA3_1 PORT MAP(
	A=> C(	3571	),
	B=>E(	3390	),
	Cin=> Carry( 	3506	),
	Cout=> Carry( 	3507	),
	S=> E(	3452	));
			
  U3508	: Soma_AMA3_1 PORT MAP(
	A=> C(	3572	),
	B=>E(	3391	),
	Cin=> Carry( 	3507	),
	Cout=> Carry( 	3508	),
	S=> E(	3453	));
			
  U3509	: Soma_AMA3_1 PORT MAP(
	A=> C(	3573	),
	B=>E(	3392	),
	Cin=> Carry( 	3508	),
	Cout=> Carry( 	3509	),
	S=> E(	3454	));
			
  U3510	: Soma_AMA3_1 PORT MAP(
	A=> C(	3574	),
	B=>E(	3393	),
	Cin=> Carry( 	3509	),
	Cout=> Carry( 	3510	),
	S=> E(	3455	));
			
  U3511	: Soma_AMA3_1 PORT MAP(
	A=> C(	3575	),
	B=>E(	3394	),
	Cin=> Carry( 	3510	),
	Cout=> Carry( 	3511	),
	S=> E(	3456	));
			
  U3512	: Soma_AMA3_1 PORT MAP(
	A=> C(	3576	),
	B=>E(	3395	),
	Cin=> Carry( 	3511	),
	Cout=> Carry( 	3512	),
	S=> E(	3457	));
			
  U3513	: Soma_AMA3_1 PORT MAP(
	A=> C(	3577	),
	B=>E(	3396	),
	Cin=> Carry( 	3512	),
	Cout=> Carry( 	3513	),
	S=> E(	3458	));
			
  U3514	: Soma_AMA3_1 PORT MAP(
	A=> C(	3578	),
	B=>E(	3397	),
	Cin=> Carry( 	3513	),
	Cout=> Carry( 	3514	),
	S=> E(	3459	));
			
  U3515	: Soma_AMA3_1 PORT MAP(
	A=> C(	3579	),
	B=>E(	3398	),
	Cin=> Carry( 	3514	),
	Cout=> Carry( 	3515	),
	S=> E(	3460	));
			
  U3516	: Soma_AMA3_1 PORT MAP(
	A=> C(	3580	),
	B=>E(	3399	),
	Cin=> Carry( 	3515	),
	Cout=> Carry( 	3516	),
	S=> E(	3461	));
			
  U3517	: Soma_AMA3_1 PORT MAP(
	A=> C(	3581	),
	B=>E(	3400	),
	Cin=> Carry( 	3516	),
	Cout=> Carry( 	3517	),
	S=> E(	3462	));
			
  U3518	: Soma_AMA3_1 PORT MAP(
	A=> C(	3582	),
	B=>E(	3401	),
	Cin=> Carry( 	3517	),
	Cout=> Carry( 	3518	),
	S=> E(	3463	));
			
  U3519	: Soma_AMA3_1 PORT MAP(
	A=> C(	3583	),
	B=>Carry(	3455	),
	Cin=> Carry( 	3518	),
	Cout=> Carry( 	3519	),
	S=> E(	3464	));

			
  U3520	: Soma_AMA3_1 PORT MAP(
	A=> C(	3584	),
	B=>E(	3402	),
	Cin=> '0'	,
	Cout=> Carry( 	3520	),
	S=> R(	56	));
			
  U3521	: Soma_AMA3_1 PORT MAP(
	A=> C(	3585	),
	B=>E(	3403	),
	Cin=> Carry( 	3520	),
	Cout=> Carry( 	3521	),
	S=> E(	3465	));
			
  U3522	: Soma_AMA3_1 PORT MAP(
	A=> C(	3586	),
	B=>E(	3404	),
	Cin=> Carry( 	3521	),
	Cout=> Carry( 	3522	),
	S=> E(	3466	));
			
  U3523	: Soma_AMA3_1 PORT MAP(
	A=> C(	3587	),
	B=>E(	3405	),
	Cin=> Carry( 	3522	),
	Cout=> Carry( 	3523	),
	S=> E(	3467	));
			
  U3524	: Soma_AMA3_1 PORT MAP(
	A=> C(	3588	),
	B=>E(	3406	),
	Cin=> Carry( 	3523	),
	Cout=> Carry( 	3524	),
	S=> E(	3468	));
			
  U3525	: Soma_AMA3_1 PORT MAP(
	A=> C(	3589	),
	B=>E(	3407	),
	Cin=> Carry( 	3524	),
	Cout=> Carry( 	3525	),
	S=> E(	3469	));
			
  U3526	: Soma_AMA3_1 PORT MAP(
	A=> C(	3590	),
	B=>E(	3408	),
	Cin=> Carry( 	3525	),
	Cout=> Carry( 	3526	),
	S=> E(	3470	));
			
  U3527	: Soma_AMA3_1 PORT MAP(
	A=> C(	3591	),
	B=>E(	3409	),
	Cin=> Carry( 	3526	),
	Cout=> Carry( 	3527	),
	S=> E(	3471	));
			
  U3528	: Soma_AMA3_1 PORT MAP(
	A=> C(	3592	),
	B=>E(	3410	),
	Cin=> Carry( 	3527	),
	Cout=> Carry( 	3528	),
	S=> E(	3472	));
			
  U3529	: Soma_AMA3_1 PORT MAP(
	A=> C(	3593	),
	B=>E(	3411	),
	Cin=> Carry( 	3528	),
	Cout=> Carry( 	3529	),
	S=> E(	3473	));
			
  U3530	: Soma_AMA3_1 PORT MAP(
	A=> C(	3594	),
	B=>E(	3412	),
	Cin=> Carry( 	3529	),
	Cout=> Carry( 	3530	),
	S=> E(	3474	));
			
  U3531	: Soma_AMA3_1 PORT MAP(
	A=> C(	3595	),
	B=>E(	3413	),
	Cin=> Carry( 	3530	),
	Cout=> Carry( 	3531	),
	S=> E(	3475	));
			
  U3532	: Soma_AMA3_1 PORT MAP(
	A=> C(	3596	),
	B=>E(	3414	),
	Cin=> Carry( 	3531	),
	Cout=> Carry( 	3532	),
	S=> E(	3476	));
			
  U3533	: Soma_AMA3_1 PORT MAP(
	A=> C(	3597	),
	B=>E(	3415	),
	Cin=> Carry( 	3532	),
	Cout=> Carry( 	3533	),
	S=> E(	3477	));
			
  U3534	: Soma_AMA3_1 PORT MAP(
	A=> C(	3598	),
	B=>E(	3416	),
	Cin=> Carry( 	3533	),
	Cout=> Carry( 	3534	),
	S=> E(	3478	));
			
  U3535	: Soma_AMA3_1 PORT MAP(
	A=> C(	3599	),
	B=>E(	3417	),
	Cin=> Carry( 	3534	),
	Cout=> Carry( 	3535	),
	S=> E(	3479	));
			
  U3536	: Soma_AMA3_1 PORT MAP(
	A=> C(	3600	),
	B=>E(	3418	),
	Cin=> Carry( 	3535	),
	Cout=> Carry( 	3536	),
	S=> E(	3480	));
			
  U3537	: Soma_AMA3_1 PORT MAP(
	A=> C(	3601	),
	B=>E(	3419	),
	Cin=> Carry( 	3536	),
	Cout=> Carry( 	3537	),
	S=> E(	3481	));
			
  U3538	: Soma_AMA3_1 PORT MAP(
	A=> C(	3602	),
	B=>E(	3420	),
	Cin=> Carry( 	3537	),
	Cout=> Carry( 	3538	),
	S=> E(	3482	));
			
  U3539	: Soma_AMA3_1 PORT MAP(
	A=> C(	3603	),
	B=>E(	3421	),
	Cin=> Carry( 	3538	),
	Cout=> Carry( 	3539	),
	S=> E(	3483	));
			
  U3540	: Soma_AMA3_1 PORT MAP(
	A=> C(	3604	),
	B=>E(	3422	),
	Cin=> Carry( 	3539	),
	Cout=> Carry( 	3540	),
	S=> E(	3484	));
			
  U3541	: Soma_AMA3_1 PORT MAP(
	A=> C(	3605	),
	B=>E(	3423	),
	Cin=> Carry( 	3540	),
	Cout=> Carry( 	3541	),
	S=> E(	3485	));
			
  U3542	: Soma_AMA3_1 PORT MAP(
	A=> C(	3606	),
	B=>E(	3424	),
	Cin=> Carry( 	3541	),
	Cout=> Carry( 	3542	),
	S=> E(	3486	));
			
  U3543	: Soma_AMA3_1 PORT MAP(
	A=> C(	3607	),
	B=>E(	3425	),
	Cin=> Carry( 	3542	),
	Cout=> Carry( 	3543	),
	S=> E(	3487	));
			
  U3544	: Soma_AMA3_1 PORT MAP(
	A=> C(	3608	),
	B=>E(	3426	),
	Cin=> Carry( 	3543	),
	Cout=> Carry( 	3544	),
	S=> E(	3488	));
			
  U3545	: Soma_AMA3_1 PORT MAP(
	A=> C(	3609	),
	B=>E(	3427	),
	Cin=> Carry( 	3544	),
	Cout=> Carry( 	3545	),
	S=> E(	3489	));
			
  U3546	: Soma_AMA3_1 PORT MAP(
	A=> C(	3610	),
	B=>E(	3428	),
	Cin=> Carry( 	3545	),
	Cout=> Carry( 	3546	),
	S=> E(	3490	));
			
  U3547	: Soma_AMA3_1 PORT MAP(
	A=> C(	3611	),
	B=>E(	3429	),
	Cin=> Carry( 	3546	),
	Cout=> Carry( 	3547	),
	S=> E(	3491	));
			
  U3548	: Soma_AMA3_1 PORT MAP(
	A=> C(	3612	),
	B=>E(	3430	),
	Cin=> Carry( 	3547	),
	Cout=> Carry( 	3548	),
	S=> E(	3492	));
			
  U3549	: Soma_AMA3_1 PORT MAP(
	A=> C(	3613	),
	B=>E(	3431	),
	Cin=> Carry( 	3548	),
	Cout=> Carry( 	3549	),
	S=> E(	3493	));
			
  U3550	: Soma_AMA3_1 PORT MAP(
	A=> C(	3614	),
	B=>E(	3432	),
	Cin=> Carry( 	3549	),
	Cout=> Carry( 	3550	),
	S=> E(	3494	));
			
  U3551	: Soma_AMA3_1 PORT MAP(
	A=> C(	3615	),
	B=>E(	3433	),
	Cin=> Carry( 	3550	),
	Cout=> Carry( 	3551	),
	S=> E(	3495	));
			
  U3552	: Soma_AMA3_1 PORT MAP(
	A=> C(	3616	),
	B=>E(	3434	),
	Cin=> Carry( 	3551	),
	Cout=> Carry( 	3552	),
	S=> E(	3496	));
			
  U3553	: Soma_AMA3_1 PORT MAP(
	A=> C(	3617	),
	B=>E(	3435	),
	Cin=> Carry( 	3552	),
	Cout=> Carry( 	3553	),
	S=> E(	3497	));
			
  U3554	: Soma_AMA3_1 PORT MAP(
	A=> C(	3618	),
	B=>E(	3436	),
	Cin=> Carry( 	3553	),
	Cout=> Carry( 	3554	),
	S=> E(	3498	));
			
  U3555	: Soma_AMA3_1 PORT MAP(
	A=> C(	3619	),
	B=>E(	3437	),
	Cin=> Carry( 	3554	),
	Cout=> Carry( 	3555	),
	S=> E(	3499	));
			
  U3556	: Soma_AMA3_1 PORT MAP(
	A=> C(	3620	),
	B=>E(	3438	),
	Cin=> Carry( 	3555	),
	Cout=> Carry( 	3556	),
	S=> E(	3500	));
			
  U3557	: Soma_AMA3_1 PORT MAP(
	A=> C(	3621	),
	B=>E(	3439	),
	Cin=> Carry( 	3556	),
	Cout=> Carry( 	3557	),
	S=> E(	3501	));
			
  U3558	: Soma_AMA3_1 PORT MAP(
	A=> C(	3622	),
	B=>E(	3440	),
	Cin=> Carry( 	3557	),
	Cout=> Carry( 	3558	),
	S=> E(	3502	));
			
  U3559	: Soma_AMA3_1 PORT MAP(
	A=> C(	3623	),
	B=>E(	3441	),
	Cin=> Carry( 	3558	),
	Cout=> Carry( 	3559	),
	S=> E(	3503	));
			
  U3560	: Soma_AMA3_1 PORT MAP(
	A=> C(	3624	),
	B=>E(	3442	),
	Cin=> Carry( 	3559	),
	Cout=> Carry( 	3560	),
	S=> E(	3504	));
			
  U3561	: Soma_AMA3_1 PORT MAP(
	A=> C(	3625	),
	B=>E(	3443	),
	Cin=> Carry( 	3560	),
	Cout=> Carry( 	3561	),
	S=> E(	3505	));
			
  U3562	: Soma_AMA3_1 PORT MAP(
	A=> C(	3626	),
	B=>E(	3444	),
	Cin=> Carry( 	3561	),
	Cout=> Carry( 	3562	),
	S=> E(	3506	));
			
  U3563	: Soma_AMA3_1 PORT MAP(
	A=> C(	3627	),
	B=>E(	3445	),
	Cin=> Carry( 	3562	),
	Cout=> Carry( 	3563	),
	S=> E(	3507	));
			
  U3564	: Soma_AMA3_1 PORT MAP(
	A=> C(	3628	),
	B=>E(	3446	),
	Cin=> Carry( 	3563	),
	Cout=> Carry( 	3564	),
	S=> E(	3508	));
			
  U3565	: Soma_AMA3_1 PORT MAP(
	A=> C(	3629	),
	B=>E(	3447	),
	Cin=> Carry( 	3564	),
	Cout=> Carry( 	3565	),
	S=> E(	3509	));
			
  U3566	: Soma_AMA3_1 PORT MAP(
	A=> C(	3630	),
	B=>E(	3448	),
	Cin=> Carry( 	3565	),
	Cout=> Carry( 	3566	),
	S=> E(	3510	));
			
  U3567	: Soma_AMA3_1 PORT MAP(
	A=> C(	3631	),
	B=>E(	3449	),
	Cin=> Carry( 	3566	),
	Cout=> Carry( 	3567	),
	S=> E(	3511	));
			
  U3568	: Soma_AMA3_1 PORT MAP(
	A=> C(	3632	),
	B=>E(	3450	),
	Cin=> Carry( 	3567	),
	Cout=> Carry( 	3568	),
	S=> E(	3512	));
			
  U3569	: Soma_AMA3_1 PORT MAP(
	A=> C(	3633	),
	B=>E(	3451	),
	Cin=> Carry( 	3568	),
	Cout=> Carry( 	3569	),
	S=> E(	3513	));
			
  U3570	: Soma_AMA3_1 PORT MAP(
	A=> C(	3634	),
	B=>E(	3452	),
	Cin=> Carry( 	3569	),
	Cout=> Carry( 	3570	),
	S=> E(	3514	));
			
  U3571	: Soma_AMA3_1 PORT MAP(
	A=> C(	3635	),
	B=>E(	3453	),
	Cin=> Carry( 	3570	),
	Cout=> Carry( 	3571	),
	S=> E(	3515	));
			
  U3572	: Soma_AMA3_1 PORT MAP(
	A=> C(	3636	),
	B=>E(	3454	),
	Cin=> Carry( 	3571	),
	Cout=> Carry( 	3572	),
	S=> E(	3516	));
			
  U3573	: Soma_AMA3_1 PORT MAP(
	A=> C(	3637	),
	B=>E(	3455	),
	Cin=> Carry( 	3572	),
	Cout=> Carry( 	3573	),
	S=> E(	3517	));
			
  U3574	: Soma_AMA3_1 PORT MAP(
	A=> C(	3638	),
	B=>E(	3456	),
	Cin=> Carry( 	3573	),
	Cout=> Carry( 	3574	),
	S=> E(	3518	));
			
  U3575	: Soma_AMA3_1 PORT MAP(
	A=> C(	3639	),
	B=>E(	3457	),
	Cin=> Carry( 	3574	),
	Cout=> Carry( 	3575	),
	S=> E(	3519	));
			
  U3576	: Soma_AMA3_1 PORT MAP(
	A=> C(	3640	),
	B=>E(	3458	),
	Cin=> Carry( 	3575	),
	Cout=> Carry( 	3576	),
	S=> E(	3520	));
			
  U3577	: Soma_AMA3_1 PORT MAP(
	A=> C(	3641	),
	B=>E(	3459	),
	Cin=> Carry( 	3576	),
	Cout=> Carry( 	3577	),
	S=> E(	3521	));
			
  U3578	: Soma_AMA3_1 PORT MAP(
	A=> C(	3642	),
	B=>E(	3460	),
	Cin=> Carry( 	3577	),
	Cout=> Carry( 	3578	),
	S=> E(	3522	));
			
  U3579	: Soma_AMA3_1 PORT MAP(
	A=> C(	3643	),
	B=>E(	3461	),
	Cin=> Carry( 	3578	),
	Cout=> Carry( 	3579	),
	S=> E(	3523	));
			
  U3580	: Soma_AMA3_1 PORT MAP(
	A=> C(	3644	),
	B=>E(	3462	),
	Cin=> Carry( 	3579	),
	Cout=> Carry( 	3580	),
	S=> E(	3524	));
			
  U3581	: Soma_AMA3_1 PORT MAP(
	A=> C(	3645	),
	B=>E(	3463	),
	Cin=> Carry( 	3580	),
	Cout=> Carry( 	3581	),
	S=> E(	3525	));
			
  U3582	: Soma_AMA3_1 PORT MAP(
	A=> C(	3646	),
	B=>E(	3464	),
	Cin=> Carry( 	3581	),
	Cout=> Carry( 	3582	),
	S=> E(	3526	));
			
  U3583	: Soma_AMA3_1 PORT MAP(
	A=> C(	3647	),
	B=>Carry(	3519	),
	Cin=> Carry( 	3582	),
	Cout=> Carry( 	3583	),
	S=> E(	3527	));

			
  U3584	: Soma_AMA3_1 PORT MAP(
	A=> C(	3648	),
	B=>E(	3465	),
	Cin=> '0'	,
	Cout=> Carry( 	3584	),
	S=> R(	57	));
			
  U3585	: Soma_AMA3_1 PORT MAP(
	A=> C(	3649	),
	B=>E(	3466	),
	Cin=> Carry( 	3584	),
	Cout=> Carry( 	3585	),
	S=> E(	3528	));
			
  U3586	: Soma_AMA3_1 PORT MAP(
	A=> C(	3650	),
	B=>E(	3467	),
	Cin=> Carry( 	3585	),
	Cout=> Carry( 	3586	),
	S=> E(	3529	));
			
  U3587	: Soma_AMA3_1 PORT MAP(
	A=> C(	3651	),
	B=>E(	3468	),
	Cin=> Carry( 	3586	),
	Cout=> Carry( 	3587	),
	S=> E(	3530	));
			
  U3588	: Soma_AMA3_1 PORT MAP(
	A=> C(	3652	),
	B=>E(	3469	),
	Cin=> Carry( 	3587	),
	Cout=> Carry( 	3588	),
	S=> E(	3531	));
			
  U3589	: Soma_AMA3_1 PORT MAP(
	A=> C(	3653	),
	B=>E(	3470	),
	Cin=> Carry( 	3588	),
	Cout=> Carry( 	3589	),
	S=> E(	3532	));
			
  U3590	: Soma_AMA3_1 PORT MAP(
	A=> C(	3654	),
	B=>E(	3471	),
	Cin=> Carry( 	3589	),
	Cout=> Carry( 	3590	),
	S=> E(	3533	));
			
  U3591	: Soma_AMA3_1 PORT MAP(
	A=> C(	3655	),
	B=>E(	3472	),
	Cin=> Carry( 	3590	),
	Cout=> Carry( 	3591	),
	S=> E(	3534	));
			
  U3592	: Soma_AMA3_1 PORT MAP(
	A=> C(	3656	),
	B=>E(	3473	),
	Cin=> Carry( 	3591	),
	Cout=> Carry( 	3592	),
	S=> E(	3535	));
			
  U3593	: Soma_AMA3_1 PORT MAP(
	A=> C(	3657	),
	B=>E(	3474	),
	Cin=> Carry( 	3592	),
	Cout=> Carry( 	3593	),
	S=> E(	3536	));
			
  U3594	: Soma_AMA3_1 PORT MAP(
	A=> C(	3658	),
	B=>E(	3475	),
	Cin=> Carry( 	3593	),
	Cout=> Carry( 	3594	),
	S=> E(	3537	));
			
  U3595	: Soma_AMA3_1 PORT MAP(
	A=> C(	3659	),
	B=>E(	3476	),
	Cin=> Carry( 	3594	),
	Cout=> Carry( 	3595	),
	S=> E(	3538	));
			
  U3596	: Soma_AMA3_1 PORT MAP(
	A=> C(	3660	),
	B=>E(	3477	),
	Cin=> Carry( 	3595	),
	Cout=> Carry( 	3596	),
	S=> E(	3539	));
			
  U3597	: Soma_AMA3_1 PORT MAP(
	A=> C(	3661	),
	B=>E(	3478	),
	Cin=> Carry( 	3596	),
	Cout=> Carry( 	3597	),
	S=> E(	3540	));
			
  U3598	: Soma_AMA3_1 PORT MAP(
	A=> C(	3662	),
	B=>E(	3479	),
	Cin=> Carry( 	3597	),
	Cout=> Carry( 	3598	),
	S=> E(	3541	));
			
  U3599	: Soma_AMA3_1 PORT MAP(
	A=> C(	3663	),
	B=>E(	3480	),
	Cin=> Carry( 	3598	),
	Cout=> Carry( 	3599	),
	S=> E(	3542	));
			
  U3600	: Soma_AMA3_1 PORT MAP(
	A=> C(	3664	),
	B=>E(	3481	),
	Cin=> Carry( 	3599	),
	Cout=> Carry( 	3600	),
	S=> E(	3543	));
			
  U3601	: Soma_AMA3_1 PORT MAP(
	A=> C(	3665	),
	B=>E(	3482	),
	Cin=> Carry( 	3600	),
	Cout=> Carry( 	3601	),
	S=> E(	3544	));
			
  U3602	: Soma_AMA3_1 PORT MAP(
	A=> C(	3666	),
	B=>E(	3483	),
	Cin=> Carry( 	3601	),
	Cout=> Carry( 	3602	),
	S=> E(	3545	));
			
  U3603	: Soma_AMA3_1 PORT MAP(
	A=> C(	3667	),
	B=>E(	3484	),
	Cin=> Carry( 	3602	),
	Cout=> Carry( 	3603	),
	S=> E(	3546	));
			
  U3604	: Soma_AMA3_1 PORT MAP(
	A=> C(	3668	),
	B=>E(	3485	),
	Cin=> Carry( 	3603	),
	Cout=> Carry( 	3604	),
	S=> E(	3547	));
			
  U3605	: Soma_AMA3_1 PORT MAP(
	A=> C(	3669	),
	B=>E(	3486	),
	Cin=> Carry( 	3604	),
	Cout=> Carry( 	3605	),
	S=> E(	3548	));
			
  U3606	: Soma_AMA3_1 PORT MAP(
	A=> C(	3670	),
	B=>E(	3487	),
	Cin=> Carry( 	3605	),
	Cout=> Carry( 	3606	),
	S=> E(	3549	));
			
  U3607	: Soma_AMA3_1 PORT MAP(
	A=> C(	3671	),
	B=>E(	3488	),
	Cin=> Carry( 	3606	),
	Cout=> Carry( 	3607	),
	S=> E(	3550	));
			
  U3608	: Soma_AMA3_1 PORT MAP(
	A=> C(	3672	),
	B=>E(	3489	),
	Cin=> Carry( 	3607	),
	Cout=> Carry( 	3608	),
	S=> E(	3551	));
			
  U3609	: Soma_AMA3_1 PORT MAP(
	A=> C(	3673	),
	B=>E(	3490	),
	Cin=> Carry( 	3608	),
	Cout=> Carry( 	3609	),
	S=> E(	3552	));
			
  U3610	: Soma_AMA3_1 PORT MAP(
	A=> C(	3674	),
	B=>E(	3491	),
	Cin=> Carry( 	3609	),
	Cout=> Carry( 	3610	),
	S=> E(	3553	));
			
  U3611	: Soma_AMA3_1 PORT MAP(
	A=> C(	3675	),
	B=>E(	3492	),
	Cin=> Carry( 	3610	),
	Cout=> Carry( 	3611	),
	S=> E(	3554	));
			
  U3612	: Soma_AMA3_1 PORT MAP(
	A=> C(	3676	),
	B=>E(	3493	),
	Cin=> Carry( 	3611	),
	Cout=> Carry( 	3612	),
	S=> E(	3555	));
			
  U3613	: Soma_AMA3_1 PORT MAP(
	A=> C(	3677	),
	B=>E(	3494	),
	Cin=> Carry( 	3612	),
	Cout=> Carry( 	3613	),
	S=> E(	3556	));
			
  U3614	: Soma_AMA3_1 PORT MAP(
	A=> C(	3678	),
	B=>E(	3495	),
	Cin=> Carry( 	3613	),
	Cout=> Carry( 	3614	),
	S=> E(	3557	));
			
  U3615	: Soma_AMA3_1 PORT MAP(
	A=> C(	3679	),
	B=>E(	3496	),
	Cin=> Carry( 	3614	),
	Cout=> Carry( 	3615	),
	S=> E(	3558	));
			
  U3616	: Soma_AMA3_1 PORT MAP(
	A=> C(	3680	),
	B=>E(	3497	),
	Cin=> Carry( 	3615	),
	Cout=> Carry( 	3616	),
	S=> E(	3559	));
			
  U3617	: Soma_AMA3_1 PORT MAP(
	A=> C(	3681	),
	B=>E(	3498	),
	Cin=> Carry( 	3616	),
	Cout=> Carry( 	3617	),
	S=> E(	3560	));
			
  U3618	: Soma_AMA3_1 PORT MAP(
	A=> C(	3682	),
	B=>E(	3499	),
	Cin=> Carry( 	3617	),
	Cout=> Carry( 	3618	),
	S=> E(	3561	));
			
  U3619	: Soma_AMA3_1 PORT MAP(
	A=> C(	3683	),
	B=>E(	3500	),
	Cin=> Carry( 	3618	),
	Cout=> Carry( 	3619	),
	S=> E(	3562	));
			
  U3620	: Soma_AMA3_1 PORT MAP(
	A=> C(	3684	),
	B=>E(	3501	),
	Cin=> Carry( 	3619	),
	Cout=> Carry( 	3620	),
	S=> E(	3563	));
			
  U3621	: Soma_AMA3_1 PORT MAP(
	A=> C(	3685	),
	B=>E(	3502	),
	Cin=> Carry( 	3620	),
	Cout=> Carry( 	3621	),
	S=> E(	3564	));
			
  U3622	: Soma_AMA3_1 PORT MAP(
	A=> C(	3686	),
	B=>E(	3503	),
	Cin=> Carry( 	3621	),
	Cout=> Carry( 	3622	),
	S=> E(	3565	));
			
  U3623	: Soma_AMA3_1 PORT MAP(
	A=> C(	3687	),
	B=>E(	3504	),
	Cin=> Carry( 	3622	),
	Cout=> Carry( 	3623	),
	S=> E(	3566	));
			
  U3624	: Soma_AMA3_1 PORT MAP(
	A=> C(	3688	),
	B=>E(	3505	),
	Cin=> Carry( 	3623	),
	Cout=> Carry( 	3624	),
	S=> E(	3567	));
			
  U3625	: Soma_AMA3_1 PORT MAP(
	A=> C(	3689	),
	B=>E(	3506	),
	Cin=> Carry( 	3624	),
	Cout=> Carry( 	3625	),
	S=> E(	3568	));
			
  U3626	: Soma_AMA3_1 PORT MAP(
	A=> C(	3690	),
	B=>E(	3507	),
	Cin=> Carry( 	3625	),
	Cout=> Carry( 	3626	),
	S=> E(	3569	));
			
  U3627	: Soma_AMA3_1 PORT MAP(
	A=> C(	3691	),
	B=>E(	3508	),
	Cin=> Carry( 	3626	),
	Cout=> Carry( 	3627	),
	S=> E(	3570	));
			
  U3628	: Soma_AMA3_1 PORT MAP(
	A=> C(	3692	),
	B=>E(	3509	),
	Cin=> Carry( 	3627	),
	Cout=> Carry( 	3628	),
	S=> E(	3571	));
			
  U3629	: Soma_AMA3_1 PORT MAP(
	A=> C(	3693	),
	B=>E(	3510	),
	Cin=> Carry( 	3628	),
	Cout=> Carry( 	3629	),
	S=> E(	3572	));
			
  U3630	: Soma_AMA3_1 PORT MAP(
	A=> C(	3694	),
	B=>E(	3511	),
	Cin=> Carry( 	3629	),
	Cout=> Carry( 	3630	),
	S=> E(	3573	));
			
  U3631	: Soma_AMA3_1 PORT MAP(
	A=> C(	3695	),
	B=>E(	3512	),
	Cin=> Carry( 	3630	),
	Cout=> Carry( 	3631	),
	S=> E(	3574	));
			
  U3632	: Soma_AMA3_1 PORT MAP(
	A=> C(	3696	),
	B=>E(	3513	),
	Cin=> Carry( 	3631	),
	Cout=> Carry( 	3632	),
	S=> E(	3575	));
			
  U3633	: Soma_AMA3_1 PORT MAP(
	A=> C(	3697	),
	B=>E(	3514	),
	Cin=> Carry( 	3632	),
	Cout=> Carry( 	3633	),
	S=> E(	3576	));
			
  U3634	: Soma_AMA3_1 PORT MAP(
	A=> C(	3698	),
	B=>E(	3515	),
	Cin=> Carry( 	3633	),
	Cout=> Carry( 	3634	),
	S=> E(	3577	));
			
  U3635	: Soma_AMA3_1 PORT MAP(
	A=> C(	3699	),
	B=>E(	3516	),
	Cin=> Carry( 	3634	),
	Cout=> Carry( 	3635	),
	S=> E(	3578	));
			
  U3636	: Soma_AMA3_1 PORT MAP(
	A=> C(	3700	),
	B=>E(	3517	),
	Cin=> Carry( 	3635	),
	Cout=> Carry( 	3636	),
	S=> E(	3579	));
			
  U3637	: Soma_AMA3_1 PORT MAP(
	A=> C(	3701	),
	B=>E(	3518	),
	Cin=> Carry( 	3636	),
	Cout=> Carry( 	3637	),
	S=> E(	3580	));
			
  U3638	: Soma_AMA3_1 PORT MAP(
	A=> C(	3702	),
	B=>E(	3519	),
	Cin=> Carry( 	3637	),
	Cout=> Carry( 	3638	),
	S=> E(	3581	));
			
  U3639	: Soma_AMA3_1 PORT MAP(
	A=> C(	3703	),
	B=>E(	3520	),
	Cin=> Carry( 	3638	),
	Cout=> Carry( 	3639	),
	S=> E(	3582	));
			
  U3640	: Soma_AMA3_1 PORT MAP(
	A=> C(	3704	),
	B=>E(	3521	),
	Cin=> Carry( 	3639	),
	Cout=> Carry( 	3640	),
	S=> E(	3583	));
			
  U3641	: Soma_AMA3_1 PORT MAP(
	A=> C(	3705	),
	B=>E(	3522	),
	Cin=> Carry( 	3640	),
	Cout=> Carry( 	3641	),
	S=> E(	3584	));
			
  U3642	: Soma_AMA3_1 PORT MAP(
	A=> C(	3706	),
	B=>E(	3523	),
	Cin=> Carry( 	3641	),
	Cout=> Carry( 	3642	),
	S=> E(	3585	));
			
  U3643	: Soma_AMA3_1 PORT MAP(
	A=> C(	3707	),
	B=>E(	3524	),
	Cin=> Carry( 	3642	),
	Cout=> Carry( 	3643	),
	S=> E(	3586	));
			
  U3644	: Soma_AMA3_1 PORT MAP(
	A=> C(	3708	),
	B=>E(	3525	),
	Cin=> Carry( 	3643	),
	Cout=> Carry( 	3644	),
	S=> E(	3587	));
			
  U3645	: Soma_AMA3_1 PORT MAP(
	A=> C(	3709	),
	B=>E(	3526	),
	Cin=> Carry( 	3644	),
	Cout=> Carry( 	3645	),
	S=> E(	3588	));
			
  U3646	: Soma_AMA3_1 PORT MAP(
	A=> C(	3710	),
	B=>E(	3527	),
	Cin=> Carry( 	3645	),
	Cout=> Carry( 	3646	),
	S=> E(	3589	));
			
  U3647	: Soma_AMA3_1 PORT MAP(
	A=> C(	3711	),
	B=>Carry(	3583	),
	Cin=> Carry( 	3646	),
	Cout=> Carry( 	3647	),
	S=> E(	3590	));


			
  U3648	: Soma_AMA3_1 PORT MAP(
	A=> C(	3712	),
	B=>E(	3528	),
	Cin=> '0'	,
	Cout=> Carry( 	3648	),
	S=> R(	58	));
			
  U3649	: Soma_AMA3_1 PORT MAP(
	A=> C(	3713	),
	B=>E(	3529	),
	Cin=> Carry( 	3648	),
	Cout=> Carry( 	3649	),
	S=> E(	3591	));
			
  U3650	: Soma_AMA3_1 PORT MAP(
	A=> C(	3714	),
	B=>E(	3530	),
	Cin=> Carry( 	3649	),
	Cout=> Carry( 	3650	),
	S=> E(	3592	));
			
  U3651	: Soma_AMA3_1 PORT MAP(
	A=> C(	3715	),
	B=>E(	3531	),
	Cin=> Carry( 	3650	),
	Cout=> Carry( 	3651	),
	S=> E(	3593	));
			
  U3652	: Soma_AMA3_1 PORT MAP(
	A=> C(	3716	),
	B=>E(	3532	),
	Cin=> Carry( 	3651	),
	Cout=> Carry( 	3652	),
	S=> E(	3594	));
			
  U3653	: Soma_AMA3_1 PORT MAP(
	A=> C(	3717	),
	B=>E(	3533	),
	Cin=> Carry( 	3652	),
	Cout=> Carry( 	3653	),
	S=> E(	3595	));
			
  U3654	: Soma_AMA3_1 PORT MAP(
	A=> C(	3718	),
	B=>E(	3534	),
	Cin=> Carry( 	3653	),
	Cout=> Carry( 	3654	),
	S=> E(	3596	));
			
  U3655	: Soma_AMA3_1 PORT MAP(
	A=> C(	3719	),
	B=>E(	3535	),
	Cin=> Carry( 	3654	),
	Cout=> Carry( 	3655	),
	S=> E(	3597	));
			
  U3656	: Soma_AMA3_1 PORT MAP(
	A=> C(	3720	),
	B=>E(	3536	),
	Cin=> Carry( 	3655	),
	Cout=> Carry( 	3656	),
	S=> E(	3598	));
			
  U3657	: Soma_AMA3_1 PORT MAP(
	A=> C(	3721	),
	B=>E(	3537	),
	Cin=> Carry( 	3656	),
	Cout=> Carry( 	3657	),
	S=> E(	3599	));
			
  U3658	: Soma_AMA3_1 PORT MAP(
	A=> C(	3722	),
	B=>E(	3538	),
	Cin=> Carry( 	3657	),
	Cout=> Carry( 	3658	),
	S=> E(	3600	));
			
  U3659	: Soma_AMA3_1 PORT MAP(
	A=> C(	3723	),
	B=>E(	3539	),
	Cin=> Carry( 	3658	),
	Cout=> Carry( 	3659	),
	S=> E(	3601	));
			
  U3660	: Soma_AMA3_1 PORT MAP(
	A=> C(	3724	),
	B=>E(	3540	),
	Cin=> Carry( 	3659	),
	Cout=> Carry( 	3660	),
	S=> E(	3602	));
			
  U3661	: Soma_AMA3_1 PORT MAP(
	A=> C(	3725	),
	B=>E(	3541	),
	Cin=> Carry( 	3660	),
	Cout=> Carry( 	3661	),
	S=> E(	3603	));
			
  U3662	: Soma_AMA3_1 PORT MAP(
	A=> C(	3726	),
	B=>E(	3542	),
	Cin=> Carry( 	3661	),
	Cout=> Carry( 	3662	),
	S=> E(	3604	));
			
  U3663	: Soma_AMA3_1 PORT MAP(
	A=> C(	3727	),
	B=>E(	3543	),
	Cin=> Carry( 	3662	),
	Cout=> Carry( 	3663	),
	S=> E(	3605	));
			
  U3664	: Soma_AMA3_1 PORT MAP(
	A=> C(	3728	),
	B=>E(	3544	),
	Cin=> Carry( 	3663	),
	Cout=> Carry( 	3664	),
	S=> E(	3606	));
			
  U3665	: Soma_AMA3_1 PORT MAP(
	A=> C(	3729	),
	B=>E(	3545	),
	Cin=> Carry( 	3664	),
	Cout=> Carry( 	3665	),
	S=> E(	3607	));
			
  U3666	: Soma_AMA3_1 PORT MAP(
	A=> C(	3730	),
	B=>E(	3546	),
	Cin=> Carry( 	3665	),
	Cout=> Carry( 	3666	),
	S=> E(	3608	));
			
  U3667	: Soma_AMA3_1 PORT MAP(
	A=> C(	3731	),
	B=>E(	3547	),
	Cin=> Carry( 	3666	),
	Cout=> Carry( 	3667	),
	S=> E(	3609	));
			
  U3668	: Soma_AMA3_1 PORT MAP(
	A=> C(	3732	),
	B=>E(	3548	),
	Cin=> Carry( 	3667	),
	Cout=> Carry( 	3668	),
	S=> E(	3610	));
			
  U3669	: Soma_AMA3_1 PORT MAP(
	A=> C(	3733	),
	B=>E(	3549	),
	Cin=> Carry( 	3668	),
	Cout=> Carry( 	3669	),
	S=> E(	3611	));
			
  U3670	: Soma_AMA3_1 PORT MAP(
	A=> C(	3734	),
	B=>E(	3550	),
	Cin=> Carry( 	3669	),
	Cout=> Carry( 	3670	),
	S=> E(	3612	));
			
  U3671	: Soma_AMA3_1 PORT MAP(
	A=> C(	3735	),
	B=>E(	3551	),
	Cin=> Carry( 	3670	),
	Cout=> Carry( 	3671	),
	S=> E(	3613	));
			
  U3672	: Soma_AMA3_1 PORT MAP(
	A=> C(	3736	),
	B=>E(	3552	),
	Cin=> Carry( 	3671	),
	Cout=> Carry( 	3672	),
	S=> E(	3614	));
			
  U3673	: Soma_AMA3_1 PORT MAP(
	A=> C(	3737	),
	B=>E(	3553	),
	Cin=> Carry( 	3672	),
	Cout=> Carry( 	3673	),
	S=> E(	3615	));
			
  U3674	: Soma_AMA3_1 PORT MAP(
	A=> C(	3738	),
	B=>E(	3554	),
	Cin=> Carry( 	3673	),
	Cout=> Carry( 	3674	),
	S=> E(	3616	));
			
  U3675	: Soma_AMA3_1 PORT MAP(
	A=> C(	3739	),
	B=>E(	3555	),
	Cin=> Carry( 	3674	),
	Cout=> Carry( 	3675	),
	S=> E(	3617	));
			
  U3676	: Soma_AMA3_1 PORT MAP(
	A=> C(	3740	),
	B=>E(	3556	),
	Cin=> Carry( 	3675	),
	Cout=> Carry( 	3676	),
	S=> E(	3618	));
			
  U3677	: Soma_AMA3_1 PORT MAP(
	A=> C(	3741	),
	B=>E(	3557	),
	Cin=> Carry( 	3676	),
	Cout=> Carry( 	3677	),
	S=> E(	3619	));
			
  U3678	: Soma_AMA3_1 PORT MAP(
	A=> C(	3742	),
	B=>E(	3558	),
	Cin=> Carry( 	3677	),
	Cout=> Carry( 	3678	),
	S=> E(	3620	));
			
  U3679	: Soma_AMA3_1 PORT MAP(
	A=> C(	3743	),
	B=>E(	3559	),
	Cin=> Carry( 	3678	),
	Cout=> Carry( 	3679	),
	S=> E(	3621	));
			
  U3680	: Soma_AMA3_1 PORT MAP(
	A=> C(	3744	),
	B=>E(	3560	),
	Cin=> Carry( 	3679	),
	Cout=> Carry( 	3680	),
	S=> E(	3622	));
			
  U3681	: Soma_AMA3_1 PORT MAP(
	A=> C(	3745	),
	B=>E(	3561	),
	Cin=> Carry( 	3680	),
	Cout=> Carry( 	3681	),
	S=> E(	3623	));
			
  U3682	: Soma_AMA3_1 PORT MAP(
	A=> C(	3746	),
	B=>E(	3562	),
	Cin=> Carry( 	3681	),
	Cout=> Carry( 	3682	),
	S=> E(	3624	));
			
  U3683	: Soma_AMA3_1 PORT MAP(
	A=> C(	3747	),
	B=>E(	3563	),
	Cin=> Carry( 	3682	),
	Cout=> Carry( 	3683	),
	S=> E(	3625	));
			
  U3684	: Soma_AMA3_1 PORT MAP(
	A=> C(	3748	),
	B=>E(	3564	),
	Cin=> Carry( 	3683	),
	Cout=> Carry( 	3684	),
	S=> E(	3626	));
			
  U3685	: Soma_AMA3_1 PORT MAP(
	A=> C(	3749	),
	B=>E(	3565	),
	Cin=> Carry( 	3684	),
	Cout=> Carry( 	3685	),
	S=> E(	3627	));
			
  U3686	: Soma_AMA3_1 PORT MAP(
	A=> C(	3750	),
	B=>E(	3566	),
	Cin=> Carry( 	3685	),
	Cout=> Carry( 	3686	),
	S=> E(	3628	));
			
  U3687	: Soma_AMA3_1 PORT MAP(
	A=> C(	3751	),
	B=>E(	3567	),
	Cin=> Carry( 	3686	),
	Cout=> Carry( 	3687	),
	S=> E(	3629	));
			
  U3688	: Soma_AMA3_1 PORT MAP(
	A=> C(	3752	),
	B=>E(	3568	),
	Cin=> Carry( 	3687	),
	Cout=> Carry( 	3688	),
	S=> E(	3630	));
			
  U3689	: Soma_AMA3_1 PORT MAP(
	A=> C(	3753	),
	B=>E(	3569	),
	Cin=> Carry( 	3688	),
	Cout=> Carry( 	3689	),
	S=> E(	3631	));
			
  U3690	: Soma_AMA3_1 PORT MAP(
	A=> C(	3754	),
	B=>E(	3570	),
	Cin=> Carry( 	3689	),
	Cout=> Carry( 	3690	),
	S=> E(	3632	));
			
  U3691	: Soma_AMA3_1 PORT MAP(
	A=> C(	3755	),
	B=>E(	3571	),
	Cin=> Carry( 	3690	),
	Cout=> Carry( 	3691	),
	S=> E(	3633	));
			
  U3692	: Soma_AMA3_1 PORT MAP(
	A=> C(	3756	),
	B=>E(	3572	),
	Cin=> Carry( 	3691	),
	Cout=> Carry( 	3692	),
	S=> E(	3634	));
			
  U3693	: Soma_AMA3_1 PORT MAP(
	A=> C(	3757	),
	B=>E(	3573	),
	Cin=> Carry( 	3692	),
	Cout=> Carry( 	3693	),
	S=> E(	3635	));
			
  U3694	: Soma_AMA3_1 PORT MAP(
	A=> C(	3758	),
	B=>E(	3574	),
	Cin=> Carry( 	3693	),
	Cout=> Carry( 	3694	),
	S=> E(	3636	));
			
  U3695	: Soma_AMA3_1 PORT MAP(
	A=> C(	3759	),
	B=>E(	3575	),
	Cin=> Carry( 	3694	),
	Cout=> Carry( 	3695	),
	S=> E(	3637	));
			
  U3696	: Soma_AMA3_1 PORT MAP(
	A=> C(	3760	),
	B=>E(	3576	),
	Cin=> Carry( 	3695	),
	Cout=> Carry( 	3696	),
	S=> E(	3638	));
			
  U3697	: Soma_AMA3_1 PORT MAP(
	A=> C(	3761	),
	B=>E(	3577	),
	Cin=> Carry( 	3696	),
	Cout=> Carry( 	3697	),
	S=> E(	3639	));
			
  U3698	: Soma_AMA3_1 PORT MAP(
	A=> C(	3762	),
	B=>E(	3578	),
	Cin=> Carry( 	3697	),
	Cout=> Carry( 	3698	),
	S=> E(	3640	));
			
  U3699	: Soma_AMA3_1 PORT MAP(
	A=> C(	3763	),
	B=>E(	3579	),
	Cin=> Carry( 	3698	),
	Cout=> Carry( 	3699	),
	S=> E(	3641	));
			
  U3700	: Soma_AMA3_1 PORT MAP(
	A=> C(	3764	),
	B=>E(	3580	),
	Cin=> Carry( 	3699	),
	Cout=> Carry( 	3700	),
	S=> E(	3642	));
			
  U3701	: Soma_AMA3_1 PORT MAP(
	A=> C(	3765	),
	B=>E(	3581	),
	Cin=> Carry( 	3700	),
	Cout=> Carry( 	3701	),
	S=> E(	3643	));
			
  U3702	: Soma_AMA3_1 PORT MAP(
	A=> C(	3766	),
	B=>E(	3582	),
	Cin=> Carry( 	3701	),
	Cout=> Carry( 	3702	),
	S=> E(	3644	));
			
  U3703	: Soma_AMA3_1 PORT MAP(
	A=> C(	3767	),
	B=>E(	3583	),
	Cin=> Carry( 	3702	),
	Cout=> Carry( 	3703	),
	S=> E(	3645	));
			
  U3704	: Soma_AMA3_1 PORT MAP(
	A=> C(	3768	),
	B=>E(	3584	),
	Cin=> Carry( 	3703	),
	Cout=> Carry( 	3704	),
	S=> E(	3646	));
			
  U3705	: Soma_AMA3_1 PORT MAP(
	A=> C(	3769	),
	B=>E(	3585	),
	Cin=> Carry( 	3704	),
	Cout=> Carry( 	3705	),
	S=> E(	3647	));
			
  U3706	: Soma_AMA3_1 PORT MAP(
	A=> C(	3770	),
	B=>E(	3586	),
	Cin=> Carry( 	3705	),
	Cout=> Carry( 	3706	),
	S=> E(	3648	));
			
  U3707	: Soma_AMA3_1 PORT MAP(
	A=> C(	3771	),
	B=>E(	3587	),
	Cin=> Carry( 	3706	),
	Cout=> Carry( 	3707	),
	S=> E(	3649	));
			
  U3708	: Soma_AMA3_1 PORT MAP(
	A=> C(	3772	),
	B=>E(	3588	),
	Cin=> Carry( 	3707	),
	Cout=> Carry( 	3708	),
	S=> E(	3650	));
			
  U3709	: Soma_AMA3_1 PORT MAP(
	A=> C(	3773	),
	B=>E(	3589	),
	Cin=> Carry( 	3708	),
	Cout=> Carry( 	3709	),
	S=> E(	3651	));
			
  U3710	: Soma_AMA3_1 PORT MAP(
	A=> C(	3774	),
	B=>E(	3590	),
	Cin=> Carry( 	3709	),
	Cout=> Carry( 	3710	),
	S=> E(	3652	));
			
  U3711	: Soma_AMA3_1 PORT MAP(
	A=> C(	3775	),
	B=>Carry(	3647	),
	Cin=> Carry( 	3710	),
	Cout=> Carry( 	3711	),
	S=> E(	3653	));

			
  U3712	: Soma_AMA3_1 PORT MAP(
	A=> C(	3776	),
	B=>E(	3591	),
	Cin=> '0'	,
	Cout=> Carry( 	3712	),
	S=> R(	59	));
			
  U3713	: Soma_AMA3_1 PORT MAP(
	A=> C(	3777	),
	B=>E(	3592	),
	Cin=> Carry( 	3712	),
	Cout=> Carry( 	3713	),
	S=> E(	3654	));
			
  U3714	: Soma_AMA3_1 PORT MAP(
	A=> C(	3778	),
	B=>E(	3593	),
	Cin=> Carry( 	3713	),
	Cout=> Carry( 	3714	),
	S=> E(	3655	));
			
  U3715	: Soma_AMA3_1 PORT MAP(
	A=> C(	3779	),
	B=>E(	3594	),
	Cin=> Carry( 	3714	),
	Cout=> Carry( 	3715	),
	S=> E(	3656	));
			
  U3716	: Soma_AMA3_1 PORT MAP(
	A=> C(	3780	),
	B=>E(	3595	),
	Cin=> Carry( 	3715	),
	Cout=> Carry( 	3716	),
	S=> E(	3657	));
			
  U3717	: Soma_AMA3_1 PORT MAP(
	A=> C(	3781	),
	B=>E(	3596	),
	Cin=> Carry( 	3716	),
	Cout=> Carry( 	3717	),
	S=> E(	3658	));
			
  U3718	: Soma_AMA3_1 PORT MAP(
	A=> C(	3782	),
	B=>E(	3597	),
	Cin=> Carry( 	3717	),
	Cout=> Carry( 	3718	),
	S=> E(	3659	));
			
  U3719	: Soma_AMA3_1 PORT MAP(
	A=> C(	3783	),
	B=>E(	3598	),
	Cin=> Carry( 	3718	),
	Cout=> Carry( 	3719	),
	S=> E(	3660	));
			
  U3720	: Soma_AMA3_1 PORT MAP(
	A=> C(	3784	),
	B=>E(	3599	),
	Cin=> Carry( 	3719	),
	Cout=> Carry( 	3720	),
	S=> E(	3661	));
			
  U3721	: Soma_AMA3_1 PORT MAP(
	A=> C(	3785	),
	B=>E(	3600	),
	Cin=> Carry( 	3720	),
	Cout=> Carry( 	3721	),
	S=> E(	3662	));
			
  U3722	: Soma_AMA3_1 PORT MAP(
	A=> C(	3786	),
	B=>E(	3601	),
	Cin=> Carry( 	3721	),
	Cout=> Carry( 	3722	),
	S=> E(	3663	));
			
  U3723	: Soma_AMA3_1 PORT MAP(
	A=> C(	3787	),
	B=>E(	3602	),
	Cin=> Carry( 	3722	),
	Cout=> Carry( 	3723	),
	S=> E(	3664	));
			
  U3724	: Soma_AMA3_1 PORT MAP(
	A=> C(	3788	),
	B=>E(	3603	),
	Cin=> Carry( 	3723	),
	Cout=> Carry( 	3724	),
	S=> E(	3665	));
			
  U3725	: Soma_AMA3_1 PORT MAP(
	A=> C(	3789	),
	B=>E(	3604	),
	Cin=> Carry( 	3724	),
	Cout=> Carry( 	3725	),
	S=> E(	3666	));
			
  U3726	: Soma_AMA3_1 PORT MAP(
	A=> C(	3790	),
	B=>E(	3605	),
	Cin=> Carry( 	3725	),
	Cout=> Carry( 	3726	),
	S=> E(	3667	));
			
  U3727	: Soma_AMA3_1 PORT MAP(
	A=> C(	3791	),
	B=>E(	3606	),
	Cin=> Carry( 	3726	),
	Cout=> Carry( 	3727	),
	S=> E(	3668	));
			
  U3728	: Soma_AMA3_1 PORT MAP(
	A=> C(	3792	),
	B=>E(	3607	),
	Cin=> Carry( 	3727	),
	Cout=> Carry( 	3728	),
	S=> E(	3669	));
			
  U3729	: Soma_AMA3_1 PORT MAP(
	A=> C(	3793	),
	B=>E(	3608	),
	Cin=> Carry( 	3728	),
	Cout=> Carry( 	3729	),
	S=> E(	3670	));
			
  U3730	: Soma_AMA3_1 PORT MAP(
	A=> C(	3794	),
	B=>E(	3609	),
	Cin=> Carry( 	3729	),
	Cout=> Carry( 	3730	),
	S=> E(	3671	));
			
  U3731	: Soma_AMA3_1 PORT MAP(
	A=> C(	3795	),
	B=>E(	3610	),
	Cin=> Carry( 	3730	),
	Cout=> Carry( 	3731	),
	S=> E(	3672	));
			
  U3732	: Soma_AMA3_1 PORT MAP(
	A=> C(	3796	),
	B=>E(	3611	),
	Cin=> Carry( 	3731	),
	Cout=> Carry( 	3732	),
	S=> E(	3673	));
			
  U3733	: Soma_AMA3_1 PORT MAP(
	A=> C(	3797	),
	B=>E(	3612	),
	Cin=> Carry( 	3732	),
	Cout=> Carry( 	3733	),
	S=> E(	3674	));
			
  U3734	: Soma_AMA3_1 PORT MAP(
	A=> C(	3798	),
	B=>E(	3613	),
	Cin=> Carry( 	3733	),
	Cout=> Carry( 	3734	),
	S=> E(	3675	));
			
  U3735	: Soma_AMA3_1 PORT MAP(
	A=> C(	3799	),
	B=>E(	3614	),
	Cin=> Carry( 	3734	),
	Cout=> Carry( 	3735	),
	S=> E(	3676	));
			
  U3736	: Soma_AMA3_1 PORT MAP(
	A=> C(	3800	),
	B=>E(	3615	),
	Cin=> Carry( 	3735	),
	Cout=> Carry( 	3736	),
	S=> E(	3677	));
			
  U3737	: Soma_AMA3_1 PORT MAP(
	A=> C(	3801	),
	B=>E(	3616	),
	Cin=> Carry( 	3736	),
	Cout=> Carry( 	3737	),
	S=> E(	3678	));
			
  U3738	: Soma_AMA3_1 PORT MAP(
	A=> C(	3802	),
	B=>E(	3617	),
	Cin=> Carry( 	3737	),
	Cout=> Carry( 	3738	),
	S=> E(	3679	));
			
  U3739	: Soma_AMA3_1 PORT MAP(
	A=> C(	3803	),
	B=>E(	3618	),
	Cin=> Carry( 	3738	),
	Cout=> Carry( 	3739	),
	S=> E(	3680	));
			
  U3740	: Soma_AMA3_1 PORT MAP(
	A=> C(	3804	),
	B=>E(	3619	),
	Cin=> Carry( 	3739	),
	Cout=> Carry( 	3740	),
	S=> E(	3681	));
			
  U3741	: Soma_AMA3_1 PORT MAP(
	A=> C(	3805	),
	B=>E(	3620	),
	Cin=> Carry( 	3740	),
	Cout=> Carry( 	3741	),
	S=> E(	3682	));
			
  U3742	: Soma_AMA3_1 PORT MAP(
	A=> C(	3806	),
	B=>E(	3621	),
	Cin=> Carry( 	3741	),
	Cout=> Carry( 	3742	),
	S=> E(	3683	));
			
  U3743	: Soma_AMA3_1 PORT MAP(
	A=> C(	3807	),
	B=>E(	3622	),
	Cin=> Carry( 	3742	),
	Cout=> Carry( 	3743	),
	S=> E(	3684	));
			
  U3744	: Soma_AMA3_1 PORT MAP(
	A=> C(	3808	),
	B=>E(	3623	),
	Cin=> Carry( 	3743	),
	Cout=> Carry( 	3744	),
	S=> E(	3685	));
			
  U3745	: Soma_AMA3_1 PORT MAP(
	A=> C(	3809	),
	B=>E(	3624	),
	Cin=> Carry( 	3744	),
	Cout=> Carry( 	3745	),
	S=> E(	3686	));
			
  U3746	: Soma_AMA3_1 PORT MAP(
	A=> C(	3810	),
	B=>E(	3625	),
	Cin=> Carry( 	3745	),
	Cout=> Carry( 	3746	),
	S=> E(	3687	));
			
  U3747	: Soma_AMA3_1 PORT MAP(
	A=> C(	3811	),
	B=>E(	3626	),
	Cin=> Carry( 	3746	),
	Cout=> Carry( 	3747	),
	S=> E(	3688	));
			
  U3748	: Soma_AMA3_1 PORT MAP(
	A=> C(	3812	),
	B=>E(	3627	),
	Cin=> Carry( 	3747	),
	Cout=> Carry( 	3748	),
	S=> E(	3689	));
			
  U3749	: Soma_AMA3_1 PORT MAP(
	A=> C(	3813	),
	B=>E(	3628	),
	Cin=> Carry( 	3748	),
	Cout=> Carry( 	3749	),
	S=> E(	3690	));
			
  U3750	: Soma_AMA3_1 PORT MAP(
	A=> C(	3814	),
	B=>E(	3629	),
	Cin=> Carry( 	3749	),
	Cout=> Carry( 	3750	),
	S=> E(	3691	));
			
  U3751	: Soma_AMA3_1 PORT MAP(
	A=> C(	3815	),
	B=>E(	3630	),
	Cin=> Carry( 	3750	),
	Cout=> Carry( 	3751	),
	S=> E(	3692	));
			
  U3752	: Soma_AMA3_1 PORT MAP(
	A=> C(	3816	),
	B=>E(	3631	),
	Cin=> Carry( 	3751	),
	Cout=> Carry( 	3752	),
	S=> E(	3693	));
			
  U3753	: Soma_AMA3_1 PORT MAP(
	A=> C(	3817	),
	B=>E(	3632	),
	Cin=> Carry( 	3752	),
	Cout=> Carry( 	3753	),
	S=> E(	3694	));
			
  U3754	: Soma_AMA3_1 PORT MAP(
	A=> C(	3818	),
	B=>E(	3633	),
	Cin=> Carry( 	3753	),
	Cout=> Carry( 	3754	),
	S=> E(	3695	));
			
  U3755	: Soma_AMA3_1 PORT MAP(
	A=> C(	3819	),
	B=>E(	3634	),
	Cin=> Carry( 	3754	),
	Cout=> Carry( 	3755	),
	S=> E(	3696	));
			
  U3756	: Soma_AMA3_1 PORT MAP(
	A=> C(	3820	),
	B=>E(	3635	),
	Cin=> Carry( 	3755	),
	Cout=> Carry( 	3756	),
	S=> E(	3697	));
			
  U3757	: Soma_AMA3_1 PORT MAP(
	A=> C(	3821	),
	B=>E(	3636	),
	Cin=> Carry( 	3756	),
	Cout=> Carry( 	3757	),
	S=> E(	3698	));
			
  U3758	: Soma_AMA3_1 PORT MAP(
	A=> C(	3822	),
	B=>E(	3637	),
	Cin=> Carry( 	3757	),
	Cout=> Carry( 	3758	),
	S=> E(	3699	));
			
  U3759	: Soma_AMA3_1 PORT MAP(
	A=> C(	3823	),
	B=>E(	3638	),
	Cin=> Carry( 	3758	),
	Cout=> Carry( 	3759	),
	S=> E(	3700	));
			
  U3760	: Soma_AMA3_1 PORT MAP(
	A=> C(	3824	),
	B=>E(	3639	),
	Cin=> Carry( 	3759	),
	Cout=> Carry( 	3760	),
	S=> E(	3701	));
			
  U3761	: Soma_AMA3_1 PORT MAP(
	A=> C(	3825	),
	B=>E(	3640	),
	Cin=> Carry( 	3760	),
	Cout=> Carry( 	3761	),
	S=> E(	3702	));
			
  U3762	: Soma_AMA3_1 PORT MAP(
	A=> C(	3826	),
	B=>E(	3641	),
	Cin=> Carry( 	3761	),
	Cout=> Carry( 	3762	),
	S=> E(	3703	));
			
  U3763	: Soma_AMA3_1 PORT MAP(
	A=> C(	3827	),
	B=>E(	3642	),
	Cin=> Carry( 	3762	),
	Cout=> Carry( 	3763	),
	S=> E(	3704	));
			
  U3764	: Soma_AMA3_1 PORT MAP(
	A=> C(	3828	),
	B=>E(	3643	),
	Cin=> Carry( 	3763	),
	Cout=> Carry( 	3764	),
	S=> E(	3705	));
			
  U3765	: Soma_AMA3_1 PORT MAP(
	A=> C(	3829	),
	B=>E(	3644	),
	Cin=> Carry( 	3764	),
	Cout=> Carry( 	3765	),
	S=> E(	3706	));
			
  U3766	: Soma_AMA3_1 PORT MAP(
	A=> C(	3830	),
	B=>E(	3645	),
	Cin=> Carry( 	3765	),
	Cout=> Carry( 	3766	),
	S=> E(	3707	));
			
  U3767	: Soma_AMA3_1 PORT MAP(
	A=> C(	3831	),
	B=>E(	3646	),
	Cin=> Carry( 	3766	),
	Cout=> Carry( 	3767	),
	S=> E(	3708	));
			
  U3768	: Soma_AMA3_1 PORT MAP(
	A=> C(	3832	),
	B=>E(	3647	),
	Cin=> Carry( 	3767	),
	Cout=> Carry( 	3768	),
	S=> E(	3709	));
			
  U3769	: Soma_AMA3_1 PORT MAP(
	A=> C(	3833	),
	B=>E(	3648	),
	Cin=> Carry( 	3768	),
	Cout=> Carry( 	3769	),
	S=> E(	3710	));
			
  U3770	: Soma_AMA3_1 PORT MAP(
	A=> C(	3834	),
	B=>E(	3649	),
	Cin=> Carry( 	3769	),
	Cout=> Carry( 	3770	),
	S=> E(	3711	));
			
  U3771	: Soma_AMA3_1 PORT MAP(
	A=> C(	3835	),
	B=>E(	3650	),
	Cin=> Carry( 	3770	),
	Cout=> Carry( 	3771	),
	S=> E(	3712	));
			
  U3772	: Soma_AMA3_1 PORT MAP(
	A=> C(	3836	),
	B=>E(	3651	),
	Cin=> Carry( 	3771	),
	Cout=> Carry( 	3772	),
	S=> E(	3713	));
			
  U3773	: Soma_AMA3_1 PORT MAP(
	A=> C(	3837	),
	B=>E(	3652	),
	Cin=> Carry( 	3772	),
	Cout=> Carry( 	3773	),
	S=> E(	3714	));
			
  U3774	: Soma_AMA3_1 PORT MAP(
	A=> C(	3838	),
	B=>E(	3653	),
	Cin=> Carry( 	3773	),
	Cout=> Carry( 	3774	),
	S=> E(	3715	));
			
  U3775	: Soma_AMA3_1 PORT MAP(
	A=> C(	3839	),
	B=>Carry(	3711	),
	Cin=> Carry( 	3774	),
	Cout=> Carry( 	3775	),
	S=> E(	3716	));


			
  U3776	: Soma_AMA3_1 PORT MAP(
	A=> C(	3840	),
	B=>E(	3654	),
	Cin=> '0'	,
	Cout=> Carry( 	3776	),
	S=> R(	60	));
			
  U3777	: Soma_AMA3_1 PORT MAP(
	A=> C(	3841	),
	B=>E(	3655	),
	Cin=> Carry( 	3776	),
	Cout=> Carry( 	3777	),
	S=> E(	3717	));
			
  U3778	: Soma_AMA3_1 PORT MAP(
	A=> C(	3842	),
	B=>E(	3656	),
	Cin=> Carry( 	3777	),
	Cout=> Carry( 	3778	),
	S=> E(	3718	));
			
  U3779	: Soma_AMA3_1 PORT MAP(
	A=> C(	3843	),
	B=>E(	3657	),
	Cin=> Carry( 	3778	),
	Cout=> Carry( 	3779	),
	S=> E(	3719	));
			
  U3780	: Soma_AMA3_1 PORT MAP(
	A=> C(	3844	),
	B=>E(	3658	),
	Cin=> Carry( 	3779	),
	Cout=> Carry( 	3780	),
	S=> E(	3720	));
			
U3781	: Soma_AMA3_1 PORT MAP(
	A=> C(	3845	),
	B=>E(	3659	),
	Cin=> Carry( 	3780	),
	Cout=> Carry( 	3781	),
	S=> E(	3721	));
			
  U3782	: Soma_AMA3_1 PORT MAP(
	A=> C(	3846	),
	B=>E(	3660	),
	Cin=> Carry( 	3781	),
	Cout=> Carry( 	3782	),
	S=> E(	3722	));
			
  U3783	: Soma_AMA3_1 PORT MAP(
	A=> C(	3847	),
	B=>E(	3661	),
	Cin=> Carry( 	3782	),
	Cout=> Carry( 	3783	),
	S=> E(	3723	));
			
  U3784	: Soma_AMA3_1 PORT MAP(
	A=> C(	3848	),
	B=>E(	3662	),
	Cin=> Carry( 	3783	),
	Cout=> Carry( 	3784	),
	S=> E(	3724	));
			
  U3785	: Soma_AMA3_1 PORT MAP(
	A=> C(	3849	),
	B=>E(	3663	),
	Cin=> Carry( 	3784	),
	Cout=> Carry( 	3785	),
	S=> E(	3725	));
			
  U3786	: Soma_AMA3_1 PORT MAP(
	A=> C(	3850	),
	B=>E(	3664	),
	Cin=> Carry( 	3785	),
	Cout=> Carry( 	3786	),
	S=> E(	3726	));
			
  U3787	: Soma_AMA3_1 PORT MAP(
	A=> C(	3851	),
	B=>E(	3665	),
	Cin=> Carry( 	3786	),
	Cout=> Carry( 	3787	),
	S=> E(	3727	));
			
  U3788	: Soma_AMA3_1 PORT MAP(
	A=> C(	3852	),
	B=>E(	3666	),
	Cin=> Carry( 	3787	),
	Cout=> Carry( 	3788	),
	S=> E(	3728	));
			
  U3789	: Soma_AMA3_1 PORT MAP(
	A=> C(	3853	),
	B=>E(	3667	),
	Cin=> Carry( 	3788	),
	Cout=> Carry( 	3789	),
	S=> E(	3729	));
			
  U3790	: Soma_AMA3_1 PORT MAP(
	A=> C(	3854	),
	B=>E(	3668	),
	Cin=> Carry( 	3789	),
	Cout=> Carry( 	3790	),
	S=> E(	3730	));
			
  U3791	: Soma_AMA3_1 PORT MAP(
	A=> C(	3855	),
	B=>E(	3669	),
	Cin=> Carry( 	3790	),
	Cout=> Carry( 	3791	),
	S=> E(	3731	));
			
  U3792	: Soma_AMA3_1 PORT MAP(
	A=> C(	3856	),
	B=>E(	3670	),
	Cin=> Carry( 	3791	),
	Cout=> Carry( 	3792	),
	S=> E(	3732	));
			
  U3793	: Soma_AMA3_1 PORT MAP(
	A=> C(	3857	),
	B=>E(	3671	),
	Cin=> Carry( 	3792	),
	Cout=> Carry( 	3793	),
	S=> E(	3733	));
			
  U3794	: Soma_AMA3_1 PORT MAP(
	A=> C(	3858	),
	B=>E(	3672	),
	Cin=> Carry( 	3793	),
	Cout=> Carry( 	3794	),
	S=> E(	3734	));
			
  U3795	: Soma_AMA3_1 PORT MAP(
	A=> C(	3859	),
	B=>E(	3673	),
	Cin=> Carry( 	3794	),
	Cout=> Carry( 	3795	),
	S=> E(	3735	));
			
  U3796	: Soma_AMA3_1 PORT MAP(
	A=> C(	3860	),
	B=>E(	3674	),
	Cin=> Carry( 	3795	),
	Cout=> Carry( 	3796	),
	S=> E(	3736	));
			
  U3797	: Soma_AMA3_1 PORT MAP(
	A=> C(	3861	),
	B=>E(	3675	),
	Cin=> Carry( 	3796	),
	Cout=> Carry( 	3797	),
	S=> E(	3737	));
			
  U3798	: Soma_AMA3_1 PORT MAP(
	A=> C(	3862	),
	B=>E(	3676	),
	Cin=> Carry( 	3797	),
	Cout=> Carry( 	3798	),
	S=> E(	3738	));
			
  U3799	: Soma_AMA3_1 PORT MAP(
	A=> C(	3863	),
	B=>E(	3677	),
	Cin=> Carry( 	3798	),
	Cout=> Carry( 	3799	),
	S=> E(	3739	));
			
  U3800	: Soma_AMA3_1 PORT MAP(
	A=> C(	3864	),
	B=>E(	3678	),
	Cin=> Carry( 	3799	),
	Cout=> Carry( 	3800	),
	S=> E(	3740	));
			
  U3801	: Soma_AMA3_1 PORT MAP(
	A=> C(	3865	),
	B=>E(	3679	),
	Cin=> Carry( 	3800	),
	Cout=> Carry( 	3801	),
	S=> E(	3741	));
			
  U3802	: Soma_AMA3_1 PORT MAP(
	A=> C(	3866	),
	B=>E(	3680	),
	Cin=> Carry( 	3801	),
	Cout=> Carry( 	3802	),
	S=> E(	3742	));
			
  U3803	: Soma_AMA3_1 PORT MAP(
	A=> C(	3867	),
	B=>E(	3681	),
	Cin=> Carry( 	3802	),
	Cout=> Carry( 	3803	),
	S=> E(	3743	));
			
  U3804	: Soma_AMA3_1 PORT MAP(
	A=> C(	3868	),
	B=>E(	3682	),
	Cin=> Carry( 	3803	),
	Cout=> Carry( 	3804	),
	S=> E(	3744	));
			
  U3805	: Soma_AMA3_1 PORT MAP(
	A=> C(	3869	),
	B=>E(	3683	),
	Cin=> Carry( 	3804	),
	Cout=> Carry( 	3805	),
	S=> E(	3745	));
			
  U3806	: Soma_AMA3_1 PORT MAP(
	A=> C(	3870	),
	B=>E(	3684	),
	Cin=> Carry( 	3805	),
	Cout=> Carry( 	3806	),
	S=> E(	3746	));
			
  U3807	: Soma_AMA3_1 PORT MAP(
	A=> C(	3871	),
	B=>E(	3685	),
	Cin=> Carry( 	3806	),
	Cout=> Carry( 	3807	),
	S=> E(	3747	));
			
  U3808	: Soma_AMA3_1 PORT MAP(
	A=> C(	3872	),
	B=>E(	3686	),
	Cin=> Carry( 	3807	),
	Cout=> Carry( 	3808	),
	S=> E(	3748	));
			
  U3809	: Soma_AMA3_1 PORT MAP(
	A=> C(	3873	),
	B=>E(	3687	),
	Cin=> Carry( 	3808	),
	Cout=> Carry( 	3809	),
	S=> E(	3749	));
			
  U3810	: Soma_AMA3_1 PORT MAP(
	A=> C(	3874	),
	B=>E(	3688	),
	Cin=> Carry( 	3809	),
	Cout=> Carry( 	3810	),
	S=> E(	3750	));
			
  U3811	: Soma_AMA3_1 PORT MAP(
	A=> C(	3875	),
	B=>E(	3689	),
	Cin=> Carry( 	3810	),
	Cout=> Carry( 	3811	),
	S=> E(	3751	));
			
  U3812	: Soma_AMA3_1 PORT MAP(
	A=> C(	3876	),
	B=>E(	3690	),
	Cin=> Carry( 	3811	),
	Cout=> Carry( 	3812	),
	S=> E(	3752	));
			
  U3813	: Soma_AMA3_1 PORT MAP(
	A=> C(	3877	),
	B=>E(	3691	),
	Cin=> Carry( 	3812	),
	Cout=> Carry( 	3813	),
	S=> E(	3753	));
			
  U3814	: Soma_AMA3_1 PORT MAP(
	A=> C(	3878	),
	B=>E(	3692	),
	Cin=> Carry( 	3813	),
	Cout=> Carry( 	3814	),
	S=> E(	3754	));
			
  U3815	: Soma_AMA3_1 PORT MAP(
	A=> C(	3879	),
	B=>E(	3693	),
	Cin=> Carry( 	3814	),
	Cout=> Carry( 	3815	),
	S=> E(	3755	));
			
  U3816	: Soma_AMA3_1 PORT MAP(
	A=> C(	3880	),
	B=>E(	3694	),
	Cin=> Carry( 	3815	),
	Cout=> Carry( 	3816	),
	S=> E(	3756	));
			
  U3817	: Soma_AMA3_1 PORT MAP(
	A=> C(	3881	),
	B=>E(	3695	),
	Cin=> Carry( 	3816	),
	Cout=> Carry( 	3817	),
	S=> E(	3757	));
			
  U3818	: Soma_AMA3_1 PORT MAP(
	A=> C(	3882	),
	B=>E(	3696	),
	Cin=> Carry( 	3817	),
	Cout=> Carry( 	3818	),
	S=> E(	3758	));
			
  U3819	: Soma_AMA3_1 PORT MAP(
	A=> C(	3883	),
	B=>E(	3697	),
	Cin=> Carry( 	3818	),
	Cout=> Carry( 	3819	),
	S=> E(	3759	));
			
  U3820	: Soma_AMA3_1 PORT MAP(
	A=> C(	3884	),
	B=>E(	3698	),
	Cin=> Carry( 	3819	),
	Cout=> Carry( 	3820	),
	S=> E(	3760	));
			
  U3821	: Soma_AMA3_1 PORT MAP(
	A=> C(	3885	),
	B=>E(	3699	),
	Cin=> Carry( 	3820	),
	Cout=> Carry( 	3821	),
	S=> E(	3761	));
			
  U3822	: Soma_AMA3_1 PORT MAP(
	A=> C(	3886	),
	B=>E(	3700	),
	Cin=> Carry( 	3821	),
	Cout=> Carry( 	3822	),
	S=> E(	3762	));
			
  U3823	: Soma_AMA3_1 PORT MAP(
	A=> C(	3887	),
	B=>E(	3701	),
	Cin=> Carry( 	3822	),
	Cout=> Carry( 	3823	),
	S=> E(	3763	));
			
  U3824	: Soma_AMA3_1 PORT MAP(
	A=> C(	3888	),
	B=>E(	3702	),
	Cin=> Carry( 	3823	),
	Cout=> Carry( 	3824	),
	S=> E(	3764	));
			
  U3825	: Soma_AMA3_1 PORT MAP(
	A=> C(	3889	),
	B=>E(	3703	),
	Cin=> Carry( 	3824	),
	Cout=> Carry( 	3825	),
	S=> E(	3765	));
			
  U3826	: Soma_AMA3_1 PORT MAP(
	A=> C(	3890	),
	B=>E(	3704	),
	Cin=> Carry( 	3825	),
	Cout=> Carry( 	3826	),
	S=> E(	3766	));
			
  U3827	: Soma_AMA3_1 PORT MAP(
	A=> C(	3891	),
	B=>E(	3705	),
	Cin=> Carry( 	3826	),
	Cout=> Carry( 	3827	),
	S=> E(	3767	));
			
  U3828	: Soma_AMA3_1 PORT MAP(
	A=> C(	3892	),
	B=>E(	3706	),
	Cin=> Carry( 	3827	),
	Cout=> Carry( 	3828	),
	S=> E(	3768	));
			
  U3829	: Soma_AMA3_1 PORT MAP(
	A=> C(	3893	),
	B=>E(	3707	),
	Cin=> Carry( 	3828	),
	Cout=> Carry( 	3829	),
	S=> E(	3769	));
			
  U3830	: Soma_AMA3_1 PORT MAP(
	A=> C(	3894	),
	B=>E(	3708	),
	Cin=> Carry( 	3829	),
	Cout=> Carry( 	3830	),
	S=> E(	3770	));
			
  U3831	: Soma_AMA3_1 PORT MAP(
	A=> C(	3895	),
	B=>E(	3709	),
	Cin=> Carry( 	3830	),
	Cout=> Carry( 	3831	),
	S=> E(	3771	));
			
  U3832	: Soma_AMA3_1 PORT MAP(
	A=> C(	3896	),
	B=>E(	3710	),
	Cin=> Carry( 	3831	),
	Cout=> Carry( 	3832	),
	S=> E(	3772	));
			
  U3833	: Soma_AMA3_1 PORT MAP(
	A=> C(	3897	),
	B=>E(	3711	),
	Cin=> Carry( 	3832	),
	Cout=> Carry( 	3833	),
	S=> E(	3773	));
			
  U3834	: Soma_AMA3_1 PORT MAP(
	A=> C(	3898	),
	B=>E(	3712	),
	Cin=> Carry( 	3833	),
	Cout=> Carry( 	3834	),
	S=> E(	3774	));
			
  U3835	: Soma_AMA3_1 PORT MAP(
	A=> C(	3899	),
	B=>E(	3713	),
	Cin=> Carry( 	3834	),
	Cout=> Carry( 	3835	),
	S=> E(	3775	));
			
  U3836	: Soma_AMA3_1 PORT MAP(
	A=> C(	3900	),
	B=>E(	3714	),
	Cin=> Carry( 	3835	),
	Cout=> Carry( 	3836	),
	S=> E(	3776	));
			
  U3837	: Soma_AMA3_1 PORT MAP(
	A=> C(	3901	),
	B=>E(	3715	),
	Cin=> Carry( 	3836	),
	Cout=> Carry( 	3837	),
	S=> E(	3777	));
			
  U3838	: Soma_AMA3_1 PORT MAP(
	A=> C(	3902	),
	B=>E(	3716	),
	Cin=> Carry( 	3837	),
	Cout=> Carry( 	3838	),
	S=> E(	3778	));
			
  U3839	: Soma_AMA3_1 PORT MAP(
	A => C(3903),
	B => Carry(3775),
	Cin => Carry(3838),
	Cout => Carry(3839),
	S => E(3779));

			
  U3840	: Soma_AMA3_1 PORT MAP(
	A=> C(	3904	),
	B=>E(	3717	),
	Cin=> '0'	,
	Cout=> Carry( 	3840	),
	S=> R(	61	));
			
  U3841	: Soma_AMA3_1 PORT MAP(
	A=> C(	3905	),
	B=>E(	3718	),
	Cin=> Carry( 	3840	),
	Cout=> Carry( 	3841	),
	S=> E(	3780	));
			
  U3842	: Soma_AMA3_1 PORT MAP(
	A=> C(	3906	),
	B=>E(	3719	),
	Cin=> Carry( 	3841	),
	Cout=> Carry( 	3842	),
	S=> E(	3781	));
			
  U3843	: Soma_AMA3_1 PORT MAP(
	A=> C(	3907	),
	B=>E(	3720	),
	Cin=> Carry( 	3842	),
	Cout=> Carry( 	3843	),
	S=> E(	3782	));
			
  U3844	: Soma_AMA3_1 PORT MAP(
	A=> C(	3908	),
	B=>E(	3721	),
	Cin=> Carry( 	3843	),
	Cout=> Carry( 	3844	),
	S=> E(	3783	));
			
  U3845	: Soma_AMA3_1 PORT MAP(
	A=> C(	3909	),
	B=>E(	3722	),
	Cin=> Carry( 	3844	),
	Cout=> Carry( 	3845	),
	S=> E(	3784	));
			
  U3846	: Soma_AMA3_1 PORT MAP(
	A=> C(	3910	),
	B=>E(	3723	),
	Cin=> Carry( 	3845	),
	Cout=> Carry( 	3846	),
	S=> E(	3785	));
			
  U3847	: Soma_AMA3_1 PORT MAP(
	A=> C(	3911	),
	B=>E(	3724	),
	Cin=> Carry( 	3846	),
	Cout=> Carry( 	3847	),
	S=> E(	3786	));
			
  U3848	: Soma_AMA3_1 PORT MAP(
	A=> C(	3912	),
	B=>E(	3725	),
	Cin=> Carry( 	3847	),
	Cout=> Carry( 	3848	),
	S=> E(	3787	));
			
  U3849	: Soma_AMA3_1 PORT MAP(
	A=> C(	3913	),
	B=>E(	3726	),
	Cin=> Carry( 	3848	),
	Cout=> Carry( 	3849	),
	S=> E(	3788	));
			
  U3850	: Soma_AMA3_1 PORT MAP(
	A=> C(	3914	),
	B=>E(	3727	),
	Cin=> Carry( 	3849	),
	Cout=> Carry( 	3850	),
	S=> E(	3789	));
			
  U3851	: Soma_AMA3_1 PORT MAP(
	A=> C(	3915	),
	B=>E(	3728	),
	Cin=> Carry( 	3850	),
	Cout=> Carry( 	3851	),
	S=> E(	3790	));
			
  U3852	: Soma_AMA3_1 PORT MAP(
	A=> C(	3916	),
	B=>E(	3729	),
	Cin=> Carry( 	3851	),
	Cout=> Carry( 	3852	),
	S=> E(	3791	));
			
  U3853	: Soma_AMA3_1 PORT MAP(
	A=> C(	3917	),
	B=>E(	3730	),
	Cin=> Carry( 	3852	),
	Cout=> Carry( 	3853	),
	S=> E(	3792	));
			
  U3854	: Soma_AMA3_1 PORT MAP(
	A=> C(	3918	),
	B=>E(	3731	),
	Cin=> Carry( 	3853	),
	Cout=> Carry( 	3854	),
	S=> E(	3793	));
			
  U3855	: Soma_AMA3_1 PORT MAP(
	A=> C(	3919	),
	B=>E(	3732	),
	Cin=> Carry( 	3854	),
	Cout=> Carry( 	3855	),
	S=> E(	3794	));
			
  U3856	: Soma_AMA3_1 PORT MAP(
	A=> C(	3920	),
	B=>E(	3733	),
	Cin=> Carry( 	3855	),
	Cout=> Carry( 	3856	),
	S=> E(	3795	));
			
  U3857	: Soma_AMA3_1 PORT MAP(
	A=> C(	3921	),
	B=>E(	3734	),
	Cin=> Carry( 	3856	),
	Cout=> Carry( 	3857	),
	S=> E(	3796	));
			
  U3858	: Soma_AMA3_1 PORT MAP(
	A=> C(	3922	),
	B=>E(	3735	),
	Cin=> Carry( 	3857	),
	Cout=> Carry( 	3858	),
	S=> E(	3797	));
			
  U3859	: Soma_AMA3_1 PORT MAP(
	A=> C(	3923	),
	B=>E(	3736	),
	Cin=> Carry( 	3858	),
	Cout=> Carry( 	3859	),
	S=> E(	3798	));
			
  U3860	: Soma_AMA3_1 PORT MAP(
	A=> C(	3924	),
	B=>E(	3737	),
	Cin=> Carry( 	3859	),
	Cout=> Carry( 	3860	),
	S=> E(	3799	));
			
  U3861	: Soma_AMA3_1 PORT MAP(
	A=> C(	3925	),
	B=>E(	3738	),
	Cin=> Carry( 	3860	),
	Cout=> Carry( 	3861	),
	S=> E(	3800	));
			
  U3862	: Soma_AMA3_1 PORT MAP(
	A=> C(	3926	),
	B=>E(	3739	),
	Cin=> Carry( 	3861	),
	Cout=> Carry( 	3862	),
	S=> E(	3801	));
			
  U3863	: Soma_AMA3_1 PORT MAP(
	A=> C(	3927	),
	B=>E(	3740	),
	Cin=> Carry( 	3862	),
	Cout=> Carry( 	3863	),
	S=> E(	3802	));
			
  U3864	: Soma_AMA3_1 PORT MAP(
	A=> C(	3928	),
	B=>E(	3741	),
	Cin=> Carry( 	3863	),
	Cout=> Carry( 	3864	),
	S=> E(	3803	));
			
  U3865	: Soma_AMA3_1 PORT MAP(
	A=> C(	3929	),
	B=>E(	3742	),
	Cin=> Carry( 	3864	),
	Cout=> Carry( 	3865	),
	S=> E(	3804	));
			
  U3866	: Soma_AMA3_1 PORT MAP(
	A=> C(	3930	),
	B=>E(	3743	),
	Cin=> Carry( 	3865	),
	Cout=> Carry( 	3866	),
	S=> E(	3805	));
			
  U3867	: Soma_AMA3_1 PORT MAP(
	A=> C(	3931	),
	B=>E(	3744	),
	Cin=> Carry( 	3866	),
	Cout=> Carry( 	3867	),
	S=> E(	3806	));
			
  U3868	: Soma_AMA3_1 PORT MAP(
	A=> C(	3932	),
	B=>E(	3745	),
	Cin=> Carry( 	3867	),
	Cout=> Carry( 	3868	),
	S=> E(	3807	));
			
  U3869	: Soma_AMA3_1 PORT MAP(
	A=> C(	3933	),
	B=>E(	3746	),
	Cin=> Carry( 	3868	),
	Cout=> Carry( 	3869	),
	S=> E(	3808	));
			
  U3870	: Soma_AMA3_1 PORT MAP(
	A=> C(	3934	),
	B=>E(	3747	),
	Cin=> Carry( 	3869	),
	Cout=> Carry( 	3870	),
	S=> E(	3809	));
			
  U3871	: Soma_AMA3_1 PORT MAP(
	A=> C(	3935	),
	B=>E(	3748	),
	Cin=> Carry( 	3870	),
	Cout=> Carry( 	3871	),
	S=> E(	3810	));
			
  U3872	: Soma_AMA3_1 PORT MAP(
	A=> C(	3936	),
	B=>E(	3749	),
	Cin=> Carry( 	3871	),
	Cout=> Carry( 	3872	),
	S=> E(	3811	));
			
  U3873	: Soma_AMA3_1 PORT MAP(
	A=> C(	3937	),
	B=>E(	3750	),
	Cin=> Carry( 	3872	),
	Cout=> Carry( 	3873	),
	S=> E(	3812	));
			
  U3874	: Soma_AMA3_1 PORT MAP(
	A=> C(	3938	),
	B=>E(	3751	),
	Cin=> Carry( 	3873	),
	Cout=> Carry( 	3874	),
	S=> E(	3813	));
			
  U3875	: Soma_AMA3_1 PORT MAP(
	A=> C(	3939	),
	B=>E(	3752	),
	Cin=> Carry( 	3874	),
	Cout=> Carry( 	3875	),
	S=> E(	3814	));
			
  U3876	: Soma_AMA3_1 PORT MAP(
	A=> C(	3940	),
	B=>E(	3753	),
	Cin=> Carry( 	3875	),
	Cout=> Carry( 	3876	),
	S=> E(	3815	));
			
  U3877	: Soma_AMA3_1 PORT MAP(
	A=> C(	3941	),
	B=>E(	3754	),
	Cin=> Carry( 	3876	),
	Cout=> Carry( 	3877	),
	S=> E(	3816	));
			
  U3878	: Soma_AMA3_1 PORT MAP(
	A=> C(	3942	),
	B=>E(	3755	),
	Cin=> Carry( 	3877	),
	Cout=> Carry( 	3878	),
	S=> E(	3817	));
			
  U3879	: Soma_AMA3_1 PORT MAP(
	A=> C(	3943	),
	B=>E(	3756	),
	Cin=> Carry( 	3878	),
	Cout=> Carry( 	3879	),
	S=> E(	3818	));
			
  U3880	: Soma_AMA3_1 PORT MAP(
	A=> C(	3944	),
	B=>E(	3757	),
	Cin=> Carry( 	3879	),
	Cout=> Carry( 	3880	),
	S=> E(	3819	));
			
  U3881	: Soma_AMA3_1 PORT MAP(
	A=> C(	3945	),
	B=>E(	3758	),
	Cin=> Carry( 	3880	),
	Cout=> Carry( 	3881	),
	S=> E(	3820	));
			
  U3882	: Soma_AMA3_1 PORT MAP(
	A=> C(	3946	),
	B=>E(	3759	),
	Cin=> Carry( 	3881	),
	Cout=> Carry( 	3882	),
	S=> E(	3821	));
			
  U3883	: Soma_AMA3_1 PORT MAP(
	A=> C(	3947	),
	B=>E(	3760	),
	Cin=> Carry( 	3882	),
	Cout=> Carry( 	3883	),
	S=> E(	3822	));
			
  U3884	: Soma_AMA3_1 PORT MAP(
	A=> C(	3948	),
	B=>E(	3761	),
	Cin=> Carry( 	3883	),
	Cout=> Carry( 	3884	),
	S=> E(	3823	));
			
  U3885	: Soma_AMA3_1 PORT MAP(
	A=> C(	3949	),
	B=>E(	3762	),
	Cin=> Carry( 	3884	),
	Cout=> Carry( 	3885	),
	S=> E(	3824	));
			
  U3886	: Soma_AMA3_1 PORT MAP(
	A=> C(	3950	),
	B=>E(	3763	),
	Cin=> Carry( 	3885	),
	Cout=> Carry( 	3886	),
	S=> E(	3825	));
			
  U3887	: Soma_AMA3_1 PORT MAP(
	A=> C(	3951	),
	B=>E(	3764	),
	Cin=> Carry( 	3886	),
	Cout=> Carry( 	3887	),
	S=> E(	3826	));
			
  U3888	: Soma_AMA3_1 PORT MAP(
	A=> C(	3952	),
	B=>E(	3765	),
	Cin=> Carry( 	3887	),
	Cout=> Carry( 	3888	),
	S=> E(	3827	));
			
  U3889	: Soma_AMA3_1 PORT MAP(
	A=> C(	3953	),
	B=>E(	3766	),
	Cin=> Carry( 	3888	),
	Cout=> Carry( 	3889	),
	S=> E(	3828	));
			
  U3890	: Soma_AMA3_1 PORT MAP(
	A=> C(	3954	),
	B=>E(	3767	),
	Cin=> Carry( 	3889	),
	Cout=> Carry( 	3890	),
	S=> E(	3829	));
			
  U3891	: Soma_AMA3_1 PORT MAP(
	A=> C(	3955	),
	B=>E(	3768	),
	Cin=> Carry( 	3890	),
	Cout=> Carry( 	3891	),
	S=> E(	3830	));
			
  U3892	: Soma_AMA3_1 PORT MAP(
	A=> C(	3956	),
	B=>E(	3769	),
	Cin=> Carry( 	3891	),
	Cout=> Carry( 	3892	),
	S=> E(	3831	));
			
  U3893	: Soma_AMA3_1 PORT MAP(
	A=> C(	3957	),
	B=>E(	3770	),
	Cin=> Carry( 	3892	),
	Cout=> Carry( 	3893	),
	S=> E(	3832	));
			
  U3894	: Soma_AMA3_1 PORT MAP(
	A=> C(	3958	),
	B=>E(	3771	),
	Cin=> Carry( 	3893	),
	Cout=> Carry( 	3894	),
	S=> E(	3833	));
			
  U3895	: Soma_AMA3_1 PORT MAP(
	A=> C(	3959	),
	B=>E(	3772	),
	Cin=> Carry( 	3894	),
	Cout=> Carry( 	3895	),
	S=> E(	3834	));
			
  U3896	: Soma_AMA3_1 PORT MAP(
	A=> C(	3960	),
	B=>E(	3773	),
	Cin=> Carry( 	3895	),
	Cout=> Carry( 	3896	),
	S=> E(	3835	));
			
  U3897	: Soma_AMA3_1 PORT MAP(
	A=> C(	3961	),
	B=>E(	3774	),
	Cin=> Carry( 	3896	),
	Cout=> Carry( 	3897	),
	S=> E(	3836	));
			
  U3898	: Soma_AMA3_1 PORT MAP(
	A=> C(	3962	),
	B=>E(	3775	),
	Cin=> Carry( 	3897	),
	Cout=> Carry( 	3898	),
	S=> E(	3837	));
			
  U3899	: Soma_AMA3_1 PORT MAP(
	A=> C(	3963	),
	B=>E(	3776	),
	Cin=> Carry( 	3898	),
	Cout=> Carry( 	3899	),
	S=> E(	3838	));
			
  U3900	: Soma_AMA3_1 PORT MAP(
	A=> C(	3964	),
	B=>E(	3777	),
	Cin=> Carry( 	3899	),
	Cout=> Carry( 	3900	),
	S=> E(	3839	));
			
  U3901	: Soma_AMA3_1 PORT MAP(
	A=> C(	3965	),
	B=>E(	3778	),
	Cin=> Carry( 	3900	),
	Cout=> Carry( 	3901	),
	S=> E(	3840	));
			
  U3902	: Soma_AMA3_1 PORT MAP(
	A=> C(	3966	),
	B=>E(	3779	),
	Cin=> Carry( 	3901	),
	Cout=> Carry( 	3902	),
	S=> E(	3841	));
			
  U3903	: Soma_AMA3_1 PORT MAP(
	A=> C(	3967	),
	B=>Carry(	3839	),
	Cin=> Carry( 	3902	),
	Cout=> Carry( 	3903	),
	S=> E(	3842	));

			
  U3904	: Soma_AMA3_1 PORT MAP(
	A=> C(	3968	),
	B=>E(	3780	),
	Cin=> '0'	,
	Cout=> Carry( 	3904	),
	S=> R(	62	));
			
  U3905	: Soma_AMA3_1 PORT MAP(
	A=> C(	3969	),
	B=>E(	3781	),
	Cin=> Carry( 	3904	),
	Cout=> Carry( 	3905	),
	S=> E(	3843	));
			
  U3906	: Soma_AMA3_1 PORT MAP(
	A=> C(	3970	),
	B=>E(	3782	),
	Cin=> Carry( 	3905	),
	Cout=> Carry( 	3906	),
	S=> E(	3844	));
			
  U3907	: Soma_AMA3_1 PORT MAP(
	A=> C(	3971	),
	B=>E(	3783	),
	Cin=> Carry( 	3906	),
	Cout=> Carry( 	3907	),
	S=> E(	3845	));
			
  U3908	: Soma_AMA3_1 PORT MAP(
	A=> C(	3972	),
	B=>E(	3784	),
	Cin=> Carry( 	3907	),
	Cout=> Carry( 	3908	),
	S=> E(	3846	));
			
  U3909	: Soma_AMA3_1 PORT MAP(
	A=> C(	3973	),
	B=>E(	3785	),
	Cin=> Carry( 	3908	),
	Cout=> Carry( 	3909	),
	S=> E(	3847	));
			
  U3910	: Soma_AMA3_1 PORT MAP(
	A=> C(	3974	),
	B=>E(	3786	),
	Cin=> Carry( 	3909	),
	Cout=> Carry( 	3910	),
	S=> E(	3848	));
			
  U3911	: Soma_AMA3_1 PORT MAP(
	A=> C(	3975	),
	B=>E(	3787	),
	Cin=> Carry( 	3910	),
	Cout=> Carry( 	3911	),
	S=> E(	3849	));
			
  U3912	: Soma_AMA3_1 PORT MAP(
	A=> C(	3976	),
	B=>E(	3788	),
	Cin=> Carry( 	3911	),
	Cout=> Carry( 	3912	),
	S=> E(	3850	));
			
  U3913	: Soma_AMA3_1 PORT MAP(
	A=> C(	3977	),
	B=>E(	3789	),
	Cin=> Carry( 	3912	),
	Cout=> Carry( 	3913	),
	S=> E(	3851	));
			
  U3914	: Soma_AMA3_1 PORT MAP(
	A=> C(	3978	),
	B=>E(	3790	),
	Cin=> Carry( 	3913	),
	Cout=> Carry( 	3914	),
	S=> E(	3852	));
			
  U3915	: Soma_AMA3_1 PORT MAP(
	A=> C(	3979	),
	B=>E(	3791	),
	Cin=> Carry( 	3914	),
	Cout=> Carry( 	3915	),
	S=> E(	3853	));
			
  U3916	: Soma_AMA3_1 PORT MAP(
	A=> C(	3980	),
	B=>E(	3792	),
	Cin=> Carry( 	3915	),
	Cout=> Carry( 	3916	),
	S=> E(	3854	));
			
  U3917	: Soma_AMA3_1 PORT MAP(
	A=> C(	3981	),
	B=>E(	3793	),
	Cin=> Carry( 	3916	),
	Cout=> Carry( 	3917	),
	S=> E(	3855	));
			
  U3918	: Soma_AMA3_1 PORT MAP(
	A=> C(	3982	),
	B=>E(	3794	),
	Cin=> Carry( 	3917	),
	Cout=> Carry( 	3918	),
	S=> E(	3856	));
			
  U3919	: Soma_AMA3_1 PORT MAP(
	A=> C(	3983	),
	B=>E(	3795	),
	Cin=> Carry( 	3918	),
	Cout=> Carry( 	3919	),
	S=> E(	3857	));
			
  U3920	: Soma_AMA3_1 PORT MAP(
	A=> C(	3984	),
	B=>E(	3796	),
	Cin=> Carry( 	3919	),
	Cout=> Carry( 	3920	),
	S=> E(	3858	));
			
  U3921	: Soma_AMA3_1 PORT MAP(
	A=> C(	3985	),
	B=>E(	3797	),
	Cin=> Carry( 	3920	),
	Cout=> Carry( 	3921	),
	S=> E(	3859	));
			
  U3922	: Soma_AMA3_1 PORT MAP(
	A=> C(	3986	),
	B=>E(	3798	),
	Cin=> Carry( 	3921	),
	Cout=> Carry( 	3922	),
	S=> E(	3860	));
			
  U3923	: Soma_AMA3_1 PORT MAP(
	A=> C(	3987	),
	B=>E(	3799	),
	Cin=> Carry( 	3922	),
	Cout=> Carry( 	3923	),
	S=> E(	3861	));
			
  U3924	: Soma_AMA3_1 PORT MAP(
	A=> C(	3988	),
	B=>E(	3800	),
	Cin=> Carry( 	3923	),
	Cout=> Carry( 	3924	),
	S=> E(	3862	));
			
  U3925	: Soma_AMA3_1 PORT MAP(
	A=> C(	3989	),
	B=>E(	3801	),
	Cin=> Carry( 	3924	),
	Cout=> Carry( 	3925	),
	S=> E(	3863	));
			
  U3926	: Soma_AMA3_1 PORT MAP(
	A=> C(	3990	),
	B=>E(	3802	),
	Cin=> Carry( 	3925	),
	Cout=> Carry( 	3926	),
	S=> E(	3864	));
			
  U3927	: Soma_AMA3_1 PORT MAP(
	A=> C(	3991	),
	B=>E(	3803	),
	Cin=> Carry( 	3926	),
	Cout=> Carry( 	3927	),
	S=> E(	3865	));
			
  U3928	: Soma_AMA3_1 PORT MAP(
	A=> C(	3992	),
	B=>E(	3804	),
	Cin=> Carry( 	3927	),
	Cout=> Carry( 	3928	),
	S=> E(	3866	));
			
  U3929	: Soma_AMA3_1 PORT MAP(
	A=> C(	3993	),
	B=>E(	3805	),
	Cin=> Carry( 	3928	),
	Cout=> Carry( 	3929	),
	S=> E(	3867	));
			
  U3930	: Soma_AMA3_1 PORT MAP(
	A=> C(	3994	),
	B=>E(	3806	),
	Cin=> Carry( 	3929	),
	Cout=> Carry( 	3930	),
	S=> E(	3868	));
			
  U3931	: Soma_AMA3_1 PORT MAP(
	A=> C(	3995	),
	B=>E(	3807	),
	Cin=> Carry( 	3930	),
	Cout=> Carry( 	3931	),
	S=> E(	3869	));
			
  U3932	: Soma_AMA3_1 PORT MAP(
	A=> C(	3996	),
	B=>E(	3808	),
	Cin=> Carry( 	3931	),
	Cout=> Carry( 	3932	),
	S=> E(	3870	));
			
  U3933	: Soma_AMA3_1 PORT MAP(
	A=> C(	3997	),
	B=>E(	3809	),
	Cin=> Carry( 	3932	),
	Cout=> Carry( 	3933	),
	S=> E(	3871	));
			
  U3934	: Soma_AMA3_1 PORT MAP(
	A=> C(	3998	),
	B=>E(	3810	),
	Cin=> Carry( 	3933	),
	Cout=> Carry( 	3934	),
	S=> E(	3872	));
			
  U3935	: Soma_AMA3_1 PORT MAP(
	A=> C(	3999	),
	B=>E(	3811	),
	Cin=> Carry( 	3934	),
	Cout=> Carry( 	3935	),
	S=> E(	3873	));
			
  U3936	: Soma_AMA3_1 PORT MAP(
	A=> C(	4000	),
	B=>E(	3812	),
	Cin=> Carry( 	3935	),
	Cout=> Carry( 	3936	),
	S=> E(	3874	));
			
  U3937	: Soma_AMA3_1 PORT MAP(
	A=> C(	4001	),
	B=>E(	3813	),
	Cin=> Carry( 	3936	),
	Cout=> Carry( 	3937	),
	S=> E(	3875	));
			
  U3938	: Soma_AMA3_1 PORT MAP(
	A=> C(	4002	),
	B=>E(	3814	),
	Cin=> Carry( 	3937	),
	Cout=> Carry( 	3938	),
	S=> E(	3876	));
			
  U3939	: Soma_AMA3_1 PORT MAP(
	A=> C(	4003	),
	B=>E(	3815	),
	Cin=> Carry( 	3938	),
	Cout=> Carry( 	3939	),
	S=> E(	3877	));
			
  U3940	: Soma_AMA3_1 PORT MAP(
	A=> C(	4004	),
	B=>E(	3816	),
	Cin=> Carry( 	3939	),
	Cout=> Carry( 	3940	),
	S=> E(	3878	));
			
  U3941	: Soma_AMA3_1 PORT MAP(
	A=> C(	4005	),
	B=>E(	3817	),
	Cin=> Carry( 	3940	),
	Cout=> Carry( 	3941	),
	S=> E(	3879	));
			
  U3942	: Soma_AMA3_1 PORT MAP(
	A=> C(	4006	),
	B=>E(	3818	),
	Cin=> Carry( 	3941	),
	Cout=> Carry( 	3942	),
	S=> E(	3880	));
			
  U3943	: Soma_AMA3_1 PORT MAP(
	A=> C(	4007	),
	B=>E(	3819	),
	Cin=> Carry( 	3942	),
	Cout=> Carry( 	3943	),
	S=> E(	3881	));
			
  U3944	: Soma_AMA3_1 PORT MAP(
	A=> C(	4008	),
	B=>E(	3820	),
	Cin=> Carry( 	3943	),
	Cout=> Carry( 	3944	),
	S=> E(	3882	));
			
  U3945	: Soma_AMA3_1 PORT MAP(
	A=> C(	4009	),
	B=>E(	3821	),
	Cin=> Carry( 	3944	),
	Cout=> Carry( 	3945	),
	S=> E(	3883	));
			
  U3946	: Soma_AMA3_1 PORT MAP(
	A=> C(	4010	),
	B=>E(	3822	),
	Cin=> Carry( 	3945	),
	Cout=> Carry( 	3946	),
	S=> E(	3884	));
			
  U3947	: Soma_AMA3_1 PORT MAP(
	A=> C(	4011	),
	B=>E(	3823	),
	Cin=> Carry( 	3946	),
	Cout=> Carry( 	3947	),
	S=> E(	3885	));
			
  U3948	: Soma_AMA3_1 PORT MAP(
	A=> C(	4012	),
	B=>E(	3824	),
	Cin=> Carry( 	3947	),
	Cout=> Carry( 	3948	),
	S=> E(	3886	));
			
  U3949	: Soma_AMA3_1 PORT MAP(
	A=> C(	4013	),
	B=>E(	3825	),
	Cin=> Carry( 	3948	),
	Cout=> Carry( 	3949	),
	S=> E(	3887	));
			
  U3950	: Soma_AMA3_1 PORT MAP(
	A=> C(	4014	),
	B=>E(	3826	),
	Cin=> Carry( 	3949	),
	Cout=> Carry( 	3950	),
	S=> E(	3888	));
			
  U3951	: Soma_AMA3_1 PORT MAP(
	A=> C(	4015	),
	B=>E(	3827	),
	Cin=> Carry( 	3950	),
	Cout=> Carry( 	3951	),
	S=> E(	3889	));
			
  U3952	: Soma_AMA3_1 PORT MAP(
	A=> C(	4016	),
	B=>E(	3828	),
	Cin=> Carry( 	3951	),
	Cout=> Carry( 	3952	),
	S=> E(	3890	));
			
  U3953	: Soma_AMA3_1 PORT MAP(
	A=> C(	4017	),
	B=>E(	3829	),
	Cin=> Carry( 	3952	),
	Cout=> Carry( 	3953	),
	S=> E(	3891	));
			
  U3954	: Soma_AMA3_1 PORT MAP(
	A=> C(	4018	),
	B=>E(	3830	),
	Cin=> Carry( 	3953	),
	Cout=> Carry( 	3954	),
	S=> E(	3892	));
			
  U3955	: Soma_AMA3_1 PORT MAP(
	A=> C(	4019	),
	B=>E(	3831	),
	Cin=> Carry( 	3954	),
	Cout=> Carry( 	3955	),
	S=> E(	3893	));
			
  U3956	: Soma_AMA3_1 PORT MAP(
	A=> C(	4020	),
	B=>E(	3832	),
	Cin=> Carry( 	3955	),
	Cout=> Carry( 	3956	),
	S=> E(	3894	));
			
  U3957	: Soma_AMA3_1 PORT MAP(
	A=> C(	4021	),
	B=>E(	3833	),
	Cin=> Carry( 	3956	),
	Cout=> Carry( 	3957	),
	S=> E(	3895	));
			
  U3958	: Soma_AMA3_1 PORT MAP(
	A=> C(	4022	),
	B=>E(	3834	),
	Cin=> Carry( 	3957	),
	Cout=> Carry( 	3958	),
	S=> E(	3896	));
 			
  U3959	: Soma_AMA3_1 PORT MAP(
	A=> C(	4023	),
	B=>E(	3835	),
	Cin=> Carry( 	3958	),
	Cout=> Carry( 	3959	),
	S=> E(	3897	));
			
  U3960	: Soma_AMA3_1 PORT MAP(
	A=> C(	4024	),
	B=>E(	3836	),
	Cin=> Carry( 	3959	),
	Cout=> Carry( 	3960	),
	S=> E(	3898	));
			
  U3961	: Soma_AMA3_1 PORT MAP(
	A=> C(	4025	),
	B=>E(	3837	),
	Cin=> Carry( 	3960	),
	Cout=> Carry( 	3961	),
	S=> E(	3899	));
			
  U3962	: Soma_AMA3_1 PORT MAP(
	A=> C(	4026	),
	B=>E(	3838	),
	Cin=> Carry( 	3961	),
	Cout=> Carry( 	3962	),
	S=> E(	3900	));
			
  U3963	: Soma_AMA3_1 PORT MAP(
	A=> C(	4027	),
	B=>E(	3839	),
	Cin=> Carry( 	3962	),
	Cout=> Carry( 	3963	),
	S=> E(	3901	));
			
  U3964	: Soma_AMA3_1 PORT MAP(
	A=> C(	4028	),
	B=>E(	3840	),
	Cin=> Carry( 	3963	),
	Cout=> Carry( 	3964	),
	S=> E(	3902	));
			
  U3965	: Soma_AMA3_1 PORT MAP(
	A=> C(	4029	),
	B=>E(	3841	),
	Cin=> Carry( 	3964	),
	Cout=> Carry( 	3965	),
	S=> E(	3903	));
			
  U3966	: Soma_AMA3_1 PORT MAP(
	A=> C(	4030	),
	B=>E(	3842	),
	Cin=> Carry( 	3965	),
	Cout=> Carry( 	3966	),
	S=> E(	3904	));
			
  U3967	: Soma_AMA3_1 PORT MAP(
	A=> C(	4031	),
	B=>Carry(	3903	),
	Cin=> Carry( 	3966	),
	Cout=> Carry( 	3967	),
	S=> E(	3905	));

			
  U3968	: Soma_AMA3_1 PORT MAP(
	A=> C(	4032	),
	B=>E(	3843	),
	Cin=> '0'	,
	Cout=> Carry( 	3968	),
	S=> R(	63	));
			
  U3969	: Soma_AMA3_1 PORT MAP(
	A=> C(	4033	),
	B=>E(	3844	),
	Cin=> Carry( 	3968	),
	Cout=> Carry( 	3969	),
	S=> R(	64	));
			
  U3970	: Soma_AMA3_1 PORT MAP(
	A=> C(	4034	),
	B=>E(	3845	),
	Cin=> Carry( 	3969	),
	Cout=> Carry( 	3970	),
	S=> R(	65	));
			
  U3971	: Soma_AMA3_1 PORT MAP(
	A=> C(	4035	),
	B=>E(	3846	),
	Cin=> Carry( 	3970	),
	Cout=> Carry( 	3971	),
	S=> R(	66	));
			
  U3972	: Soma_AMA3_1 PORT MAP(
	A=> C(	4036	),
	B=>E(	3847	),
	Cin=> Carry( 	3971	),
	Cout=> Carry( 	3972	),
	S=> R(	67	));
			
  U3973	: Soma_AMA3_1 PORT MAP(
	A=> C(	4037	),
	B=>E(	3848	),
	Cin=> Carry( 	3972	),
	Cout=> Carry( 	3973	),
	S=> R(	68	));
			
  U3974	: Soma_AMA3_1 PORT MAP(
	A=> C(	4038	),
	B=>E(	3849	),
	Cin=> Carry( 	3973	),
	Cout=> Carry( 	3974	),
	S=> R(	69	));
			
  U3975	: Soma_AMA3_1 PORT MAP(
	A=> C(	4039	),
	B=>E(	3850	),
	Cin=> Carry( 	3974	),
	Cout=> Carry( 	3975	),
	S=> R(	70	));
			
  U3976	: Soma_AMA3_1 PORT MAP(
	A=> C(	4040	),
	B=>E(	3851	),
	Cin=> Carry( 	3975	),
	Cout=> Carry( 	3976	),
	S=> R(	71	));
			
  U3977	: Soma_AMA3_1 PORT MAP(
	A=> C(	4041	),
	B=>E(	3852	),
	Cin=> Carry( 	3976	),
	Cout=> Carry( 	3977	),
	S=> R(	72	));
			
  U3978	: Soma_AMA3_1 PORT MAP(
	A=> C(	4042	),
	B=>E(	3853	),
	Cin=> Carry( 	3977	),
	Cout=> Carry( 	3978	),
	S=> R(	73	));
			
  U3979	: Soma_AMA3_1 PORT MAP(
	A=> C(	4043	),
	B=>E(	3854	),
	Cin=> Carry( 	3978	),
	Cout=> Carry( 	3979	),
	S=> R(	74	));
			
  U3980	: Soma_AMA3_1 PORT MAP(
	A=> C(	4044	),
	B=>E(	3855	),
	Cin=> Carry( 	3979	),
	Cout=> Carry( 	3980	),
	S=> R(	75	));
			
  U3981	: Soma_AMA3_1 PORT MAP(
	A=> C(	4045	),
	B=>E(	3856	),
	Cin=> Carry( 	3980	),
	Cout=> Carry( 	3981	),
	S=> R(	76	));
			
  U3982	: Soma_AMA3_1 PORT MAP(
	A=> C(	4046	),
	B=>E(	3857	),
	Cin=> Carry( 	3981	),
	Cout=> Carry( 	3982	),
	S=> R(	77	));
			
  U3983	: Soma_AMA3_1 PORT MAP(
	A=> C(	4047	),
	B=>E(	3858	),
	Cin=> Carry( 	3982	),
	Cout=> Carry( 	3983	),
	S=> R(	78	));
			
  U3984	: Soma_AMA3_1 PORT MAP(
	A=> C(	4048	),
	B=>E(	3859	),
	Cin=> Carry( 	3983	),
	Cout=> Carry( 	3984	),
	S=> R(	79	));
			
  U3985	: Soma_AMA3_1 PORT MAP(
	A=> C(	4049	),
	B=>E(	3860	),
	Cin=> Carry( 	3984	),
	Cout=> Carry( 	3985	),
	S=> R(	80	));
			
  U3986	: Soma_AMA3_1 PORT MAP(
	A=> C(	4050	),
	B=>E(	3861	),
	Cin=> Carry( 	3985	),
	Cout=> Carry( 	3986	),
	S=> R(	81	));
			
  U3987	: Soma_AMA3_1 PORT MAP(
	A=> C(	4051	),
	B=>E(	3862	),
	Cin=> Carry( 	3986	),
	Cout=> Carry( 	3987	),
	S=> R(	82	));
			
  U3988	: Soma_AMA3_1 PORT MAP(
	A=> C(	4052	),
	B=>E(	3863	),
	Cin=> Carry( 	3987	),
	Cout=> Carry( 	3988	),
	S=> R(	83	));
			
  U3989	: Soma_AMA3_1 PORT MAP(
	A=> C(	4053	),
	B=>E(	3864	),
	Cin=> Carry( 	3988	),
	Cout=> Carry( 	3989	),
	S=> R(	84	));
			
  U3990	: Soma_AMA3_1 PORT MAP(
	A=> C(	4054	),
	B=>E(	3865	),
	Cin=> Carry( 	3989	),
	Cout=> Carry( 	3990	),
	S=> R(	85	));
			
  U3991	: Soma_AMA3_1 PORT MAP(
	A=> C(	4055	),
	B=>E(	3866	),
	Cin=> Carry( 	3990	),
	Cout=> Carry( 	3991	),
	S=> R(	86	));
			
  U3992	: Soma_AMA3_1 PORT MAP(
	A=> C(	4056	),
	B=>E(	3867	),
	Cin=> Carry( 	3991	),
	Cout=> Carry( 	3992	),
	S=> R(	87	));
			
  U3993	: Soma_AMA3_1 PORT MAP(
	A=> C(	4057	),
	B=>E(	3868	),
	Cin=> Carry( 	3992	),
	Cout=> Carry( 	3993	),
	S=> R(	88	));
			
  U3994	: Soma_AMA3_1 PORT MAP(
	A=> C(	4058	),
	B=>E(	3869	),
	Cin=> Carry( 	3993	),
	Cout=> Carry( 	3994	),
	S=> R(	89	));
			
  U3995	: Soma_AMA3_1 PORT MAP(
	A=> C(	4059	),
	B=>E(	3870	),
	Cin=> Carry( 	3994	),
	Cout=> Carry( 	3995	),
	S=> R(	90	));
			
  U3996	: Soma_AMA3_1 PORT MAP(
	A=> C(	4060	),
	B=>E(	3871	),
	Cin=> Carry( 	3995	),
	Cout=> Carry( 	3996	),
	S=> R(	91	));
			
  U3997	: Soma_AMA3_1 PORT MAP(
	A=> C(	4061	),
	B=>E(	3872	),
	Cin=> Carry( 	3996	),
	Cout=> Carry( 	3997	),
	S=> R(	92	));
			
  U3998	: Soma_AMA3_1 PORT MAP(
	A=> C(	4062	),
	B=>E(	3873	),
	Cin=> Carry( 	3997	),
	Cout=> Carry( 	3998	),
	S=> R(	93	));
			
  U3999	: Soma_AMA3_1 PORT MAP(
	A=> C(	4063	),
	B=>E(	3874	),
	Cin=> Carry( 	3998	),
	Cout=> Carry( 	3999	),
	S=> R(	94	));
			
  U4000	: Soma_AMA3_1 PORT MAP(
	A=> C(	4064	),
	B=>E(	3875	),
	Cin=> Carry( 	3999	),
	Cout=> Carry( 	4000	),
	S=> R(	95	));
			
  U4001	: Soma_AMA3_1 PORT MAP(
	A=> C(	4065	),
	B=>E(	3876	),
	Cin=> Carry( 	4000	),
	Cout=> Carry( 	4001	),
	S=> R(	96	));
			
  U4002	: Soma_AMA3_1 PORT MAP(
	A=> C(	4066	),
	B=>E(	3877	),
	Cin=> Carry( 	4001	),
	Cout=> Carry( 	4002	),
	S=> R(	97	));
			
  U4003	: Soma_AMA3_1 PORT MAP(
	A=> C(	4067	),
	B=>E(	3878	),
	Cin=> Carry( 	4002	),
	Cout=> Carry( 	4003	),
	S=> R(	98	));
			
  U4004	: Soma_AMA3_1 PORT MAP(
	A=> C(	4068	),
	B=>E(	3879	),
	Cin=> Carry( 	4003	),
	Cout=> Carry( 	4004	),
	S=> R(	99	));
			
  U4005	: Soma_AMA3_1 PORT MAP(
	A=> C(	4069	),
	B=>E(	3880	),
	Cin=> Carry( 	4004	),
	Cout=> Carry( 	4005	),
	S=> R(	100	));
			
  U4006	: Soma_AMA3_1 PORT MAP(
	A=> C(	4070	),
	B=>E(	3881	),
	Cin=> Carry( 	4005	),
	Cout=> Carry( 	4006	),
	S=> R(	101	));
			
  U4007	: Soma_AMA3_1 PORT MAP(
	A=> C(	4071	),
	B=>E(	3882	),
	Cin=> Carry( 	4006	),
	Cout=> Carry( 	4007	),
	S=> R(	102	));
			
  U4008	: Soma_AMA3_1 PORT MAP(
	A=> C(	4072	),
	B=>E(	3883	),
	Cin=> Carry( 	4007	),
	Cout=> Carry( 	4008	),
	S=> R(	103	));
			
  U4009	: Soma_AMA3_1 PORT MAP(
	A=> C(	4073	),
	B=>E(	3884	),
	Cin=> Carry( 	4008	),
	Cout=> Carry( 	4009	),
	S=> R(	104	));
			
  U4010	: Soma_AMA3_1 PORT MAP(
	A=> C(	4074	),
	B=>E(	3885	),
	Cin=> Carry( 	4009	),
	Cout=> Carry( 	4010	),
	S=> R(	105	));
			
  U4011	: Soma_AMA3_1 PORT MAP(
	A=> C(	4075	),
	B=>E(	3886	),
	Cin=> Carry( 	4010	),
	Cout=> Carry( 	4011	),
	S=> R(	106	));
			
  U4012	: Soma_AMA3_1 PORT MAP(
	A=> C(	4076	),
	B=>E(	3887	),
	Cin=> Carry( 	4011	),
	Cout=> Carry( 	4012	),
	S=> R(	107	));
			
  U4013	: Soma_AMA3_1 PORT MAP(
	A=> C(	4077	),
	B=>E(	3888	),
	Cin=> Carry( 	4012	),
	Cout=> Carry( 	4013	),
	S=> R(	108	));
			
  U4014	: Soma_AMA3_1 PORT MAP(
	A=> C(	4078	),
	B=>E(	3889	),
	Cin=> Carry( 	4013	),
	Cout=> Carry( 	4014	),
	S=> R(	109	));
			
  U4015	: Soma_AMA3_1 PORT MAP(
	A=> C(	4079	),
	B=>E(	3890	),
	Cin=> Carry( 	4014	),
	Cout=> Carry( 	4015	),
	S=> R(	110	));
			
  U4016	: Soma_AMA3_1 PORT MAP(
	A=> C(	4080	),
	B=>E(	3891	),
	Cin=> Carry( 	4015	),
	Cout=> Carry( 	4016	),
	S=> R(	111	));
			
  U4017	: Soma_AMA3_1 PORT MAP(
	A=> C(	4081	),
	B=>E(	3892	),
	Cin=> Carry( 	4016	),
	Cout=> Carry( 	4017	),
	S=> R(	112	));
			
  U4018	: Soma_AMA3_1 PORT MAP(
	A=> C(	4082	),
	B=>E(	3893	),
	Cin=> Carry( 	4017	),
	Cout=> Carry( 	4018	),
	S=> R(	113	));
			
  U4019	: Soma_AMA3_1 PORT MAP(
	A=> C(	4083	),
	B=>E(	3894	),
	Cin=> Carry( 	4018	),
	Cout=> Carry( 	4019	),
	S=> R(	114	));
			
  U4020	: Soma_AMA3_1 PORT MAP(
	A=> C(	4084	),
	B=>E(	3895	),
	Cin=> Carry( 	4019	),
	Cout=> Carry( 	4020	),
	S=> R(	115	));
			
  U4021	: Soma_AMA3_1 PORT MAP(
	A=> C(	4085	),
	B=>E(	3896	),
	Cin=> Carry( 	4020	),
	Cout=> Carry( 	4021	),
	S=> R(	116	));
			
  U4022	: Soma_AMA3_1 PORT MAP(
	A=> C(	4086	),
	B=>E(	3897	),
	Cin=> Carry( 	4021	),
	Cout=> Carry( 	4022	),
	S=> R(	117	));
			
  U4023	: Soma_AMA3_1 PORT MAP(
	A=> C(	4087	),
	B=>E(	3898	),
	Cin=> Carry( 	4022	),
	Cout=> Carry( 	4023	),
	S=> R(	118	));
			
  U4024	: Soma_AMA3_1 PORT MAP(
	A=> C(	4088	),
	B=>E(	3899	),
	Cin=> Carry( 	4023	),
	Cout=> Carry( 	4024	),
	S=> R(	119	));
			
  U4025	: Soma_AMA3_1 PORT MAP(
	A=> C(	4089	),
	B=>E(	3900	),
	Cin=> Carry( 	4024	),
	Cout=> Carry( 	4025	),
	S=> R(	120	));
			
  U4026	: Soma_AMA3_1 PORT MAP(
	A=> C(	4090	),
	B=>E(	3901	),
	Cin=> Carry( 	4025	),
	Cout=> Carry( 	4026	),
	S=> R(	121	));
			
  U4027	: Soma_AMA3_1 PORT MAP(
	A=> C(	4091	),
	B=>E(	3902	),
	Cin=> Carry( 	4026	),
	Cout=> Carry( 	4027	),
	S=> R(	122	));
			
  U4028	: Soma_AMA3_1 PORT MAP(
	A=> C(	4092	),
	B=>E(	3903	),
	Cin=> Carry( 	4027	),
	Cout=> Carry( 	4028	),
	S=> R(	123	));
			
  U4029	: Soma_AMA3_1 PORT MAP(
	A=> C(	4093	),
	B=>E(	3904	),
	Cin=> Carry( 	4028	),
	Cout=> Carry( 	4029	),
	S=> R(	124	));
			
  U4030	: Soma_AMA3_1 PORT MAP(
	A=> C(	4094	),
	B=>E(	3905	),
	Cin=> Carry( 	4029	),
	Cout=> Carry( 	4030	),
	S=> R(	125	));
			
  U4031	: Soma_AMA3_1 PORT MAP(
	A => C(4095),
	B => Carry(3967),
	Cin => Carry(4030),
	Cout => R(127),
	S => R(126));





  
end Mult64;

